
module ddr2_init_engine_DW01_inc_1 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n5, n6, n9, n12, n13, n14, n17, n18, n21, n22, n25, n28, n29, n30,
         n31, n34, n37, n38, n39, n40, n41, n42, n43, n44;

  NAND2X1 U5 ( .A(A[0]), .B(A[1]), .Y(n5) );
  NAND2X1 U10 ( .A(A[2]), .B(n6), .Y(n9) );
  NAND2X1 U14 ( .A(A[3]), .B(A[2]), .Y(n12) );
  NOR2X1 U15 ( .A(n5), .B(n12), .Y(n13) );
  NOR2X1 U21 ( .A(n17), .B(n14), .Y(n18) );
  XOR2X1 U22 ( .A(n14), .B(n17), .Y(SUM[4]) );
  NAND2X1 U25 ( .A(A[4]), .B(A[5]), .Y(n21) );
  NOR2X1 U26 ( .A(n21), .B(n14), .Y(n22) );
  NAND2X1 U30 ( .A(A[6]), .B(n22), .Y(n25) );
  NAND2X1 U34 ( .A(A[6]), .B(A[7]), .Y(n28) );
  NOR2X1 U35 ( .A(n21), .B(n28), .Y(n29) );
  NAND2X1 U36 ( .A(n13), .B(n29), .Y(n30) );
  NAND2X1 U41 ( .A(A[8]), .B(n31), .Y(n34) );
  NAND2X1 U45 ( .A(A[9]), .B(A[8]), .Y(n37) );
  NOR2X1 U46 ( .A(n37), .B(n30), .Y(n38) );
  HAX1 U48 ( .A(A[10]), .B(n38), .YC(n39), .YS(SUM[10]) );
  HAX1 U49 ( .A(A[11]), .B(n39), .YC(n40), .YS(SUM[11]) );
  HAX1 U50 ( .A(A[12]), .B(n40), .YC(n41), .YS(SUM[12]) );
  HAX1 U51 ( .A(A[13]), .B(n41), .YC(n42), .YS(SUM[13]) );
  HAX1 U52 ( .A(A[14]), .B(n42), .YC(n43), .YS(SUM[14]) );
  HAX1 U53 ( .A(A[15]), .B(n43), .YC(n44), .YS(SUM[15]) );
  XOR2X1 U54 ( .A(n44), .B(A[16]), .Y(SUM[16]) );
  XNOR2X1 U57 ( .A(n9), .B(A[3]), .Y(SUM[3]) );
  XOR2X1 U58 ( .A(A[2]), .B(n6), .Y(SUM[2]) );
  XOR2X1 U59 ( .A(A[1]), .B(A[0]), .Y(SUM[1]) );
  XOR2X1 U60 ( .A(n18), .B(A[5]), .Y(SUM[5]) );
  XOR2X1 U61 ( .A(n22), .B(A[6]), .Y(SUM[6]) );
  XNOR2X1 U62 ( .A(n25), .B(A[7]), .Y(SUM[7]) );
  XOR2X1 U63 ( .A(n31), .B(A[8]), .Y(SUM[8]) );
  XNOR2X1 U64 ( .A(n34), .B(A[9]), .Y(SUM[9]) );
  INVX2 U65 ( .A(n5), .Y(n6) );
  INVX2 U66 ( .A(n30), .Y(n31) );
  INVX2 U67 ( .A(A[4]), .Y(n17) );
  INVX2 U68 ( .A(n13), .Y(n14) );
  INVX2 U69 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DEPTH_P26_WIDTH16_DW01_inc_2 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   carry_5_, carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_4 ( .A(A[4]), .B(carry_4_), .YC(carry_5_), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry_5_), .B(A[5]), .Y(SUM[5]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DEPTH_P26_WIDTH16_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;
  wire   carry_6_, carry_5_, carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_5 ( .A(A[5]), .B(carry_5_), .YC(carry_6_), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry_4_), .YC(carry_5_), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry_6_), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DEPTH_P26_WIDTH16_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   carry_5_, carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_4 ( .A(A[4]), .B(carry_4_), .YC(carry_5_), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry_5_), .B(A[5]), .Y(SUM[5]) );
endmodule


module FIFO_DEPTH_P26_WIDTH16_DW01_dec_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  XOR2X1 U1 ( .A(A[6]), .B(n1), .Y(SUM[6]) );
  NOR2X1 U2 ( .A(A[5]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[5]), .B(n2), .Y(SUM[5]) );
  OAI21X1 U4 ( .A(n3), .B(n4), .C(n2), .Y(SUM[4]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[4]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[3]) );
  AOI21X1 U8 ( .A(n6), .B(A[3]), .C(n3), .Y(n5) );
  NOR2X1 U9 ( .A(n6), .B(A[3]), .Y(n3) );
  OAI21X1 U10 ( .A(n7), .B(n8), .C(n6), .Y(SUM[2]) );
  NAND2X1 U11 ( .A(n7), .B(n8), .Y(n6) );
  INVX1 U12 ( .A(A[2]), .Y(n8) );
  INVX1 U13 ( .A(n9), .Y(SUM[1]) );
  AOI21X1 U14 ( .A(A[0]), .B(A[1]), .C(n7), .Y(n9) );
  NOR2X1 U15 ( .A(A[1]), .B(A[0]), .Y(n7) );
  INVX1 U16 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DEPTH_P26_WIDTH33_DW01_inc_2 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   carry_5_, carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_4 ( .A(A[4]), .B(carry_4_), .YC(carry_5_), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry_5_), .B(A[5]), .Y(SUM[5]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DEPTH_P26_WIDTH33_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;
  wire   carry_6_, carry_5_, carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_5 ( .A(A[5]), .B(carry_5_), .YC(carry_6_), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry_4_), .YC(carry_5_), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry_6_), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DEPTH_P26_WIDTH33_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   carry_5_, carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_4 ( .A(A[4]), .B(carry_4_), .YC(carry_5_), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry_5_), .B(A[5]), .Y(SUM[5]) );
endmodule


module FIFO_DEPTH_P26_WIDTH33_DW01_dec_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  XOR2X1 U1 ( .A(A[6]), .B(n1), .Y(SUM[6]) );
  NOR2X1 U2 ( .A(A[5]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[5]), .B(n2), .Y(SUM[5]) );
  OAI21X1 U4 ( .A(n3), .B(n4), .C(n2), .Y(SUM[4]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[4]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[3]) );
  AOI21X1 U8 ( .A(n6), .B(A[3]), .C(n3), .Y(n5) );
  NOR2X1 U9 ( .A(n6), .B(A[3]), .Y(n3) );
  OAI21X1 U10 ( .A(n7), .B(n8), .C(n6), .Y(SUM[2]) );
  NAND2X1 U11 ( .A(n7), .B(n8), .Y(n6) );
  INVX1 U12 ( .A(A[2]), .Y(n8) );
  INVX1 U13 ( .A(n9), .Y(SUM[1]) );
  AOI21X1 U14 ( .A(A[0]), .B(A[1]), .C(n7), .Y(n9) );
  NOR2X1 U15 ( .A(A[1]), .B(A[0]), .Y(n7) );
  INVX1 U16 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DEPTH_P26_WIDTH41_DW01_inc_2 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   carry_5_, carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_4 ( .A(A[4]), .B(carry_4_), .YC(carry_5_), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry_5_), .B(A[5]), .Y(SUM[5]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DEPTH_P26_WIDTH41_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;
  wire   carry_6_, carry_5_, carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_5 ( .A(A[5]), .B(carry_5_), .YC(carry_6_), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry_4_), .YC(carry_5_), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry_6_), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIFO_DEPTH_P26_WIDTH41_DW01_inc_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   carry_5_, carry_4_, carry_3_, carry_2_;

  HAX1 U1_1_4 ( .A(A[4]), .B(carry_4_), .YC(carry_5_), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry_3_), .YC(carry_4_), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry_2_), .YC(carry_3_), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry_2_), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry_5_), .B(A[5]), .Y(SUM[5]) );
endmodule


module FIFO_DEPTH_P26_WIDTH41_DW01_dec_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  XOR2X1 U1 ( .A(A[6]), .B(n1), .Y(SUM[6]) );
  NOR2X1 U2 ( .A(A[5]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[5]), .B(n2), .Y(SUM[5]) );
  OAI21X1 U4 ( .A(n3), .B(n4), .C(n2), .Y(SUM[4]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[4]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[3]) );
  AOI21X1 U8 ( .A(n6), .B(A[3]), .C(n3), .Y(n5) );
  NOR2X1 U9 ( .A(n6), .B(A[3]), .Y(n3) );
  OAI21X1 U10 ( .A(n7), .B(n8), .C(n6), .Y(SUM[2]) );
  NAND2X1 U11 ( .A(n7), .B(n8), .Y(n6) );
  INVX1 U12 ( .A(A[2]), .Y(n8) );
  INVX1 U13 ( .A(n9), .Y(SUM[1]) );
  AOI21X1 U14 ( .A(A[0]), .B(A[1]), .C(n7), .Y(n9) );
  NOR2X1 U15 ( .A(A[1]), .B(A[0]), .Y(n7) );
  INVX1 U16 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SSTL18DDR2_41 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_40 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_39 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_38 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_37 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_36 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_35 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_34 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_33 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_32 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_31 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_30 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_29 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_28 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_27 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_26 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_25 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_24 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_23 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_22 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_21 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_20 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_19 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_18 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_17 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_16 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_15 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_14 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_13 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_12 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_11 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_10 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_9 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_8 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_7 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_6 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_5 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_4 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_3 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_2 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_1 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_0 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX1 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR2_42 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX1 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
  INVX2 U1 ( .A(A), .Y(n2) );
endmodule


module SSTL18DDR2DIFF ( PAD, PADN, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD,  PADN;
  wire   n4, n5, n6;

  TBUFX1 b2 ( .A(A), .EN(TS), .Y(PADN) );
  TBUFX1 b1 ( .A(n6), .EN(TS), .Y(PAD) );
  NAND3X1 U3 ( .A(PAD), .B(n5), .C(RI), .Y(n4) );
  INVX2 U1 ( .A(A), .Y(n6) );
  INVX2 U2 ( .A(n4), .Y(Z) );
  INVX2 U4 ( .A(PADN), .Y(n5) );
endmodule


module SSTL18DDR2INTERFACE ( ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, 
        casbar_pad, webar_pad, ba_pad, a_pad, dm_pad, odt_pad, dq_o, dqs_o, 
        dqsbar_o, dq_pad, dqs_pad, dqsbar_pad, ri_i, ts_i, ck_i, cke_i, 
        csbar_i, rasbar_i, casbar_i, webar_i, ba_i, a_i, dq_i, dqs_i, dqsbar_i, 
        dm_i, odt_i );
  output [1:0] ba_pad;
  output [12:0] a_pad;
  output [1:0] dm_pad;
  output [15:0] dq_o;
  output [1:0] dqs_o;
  output [1:0] dqsbar_o;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [1:0] ba_i;
  input [12:0] a_i;
  input [15:0] dq_i;
  input [1:0] dqs_i;
  input [1:0] dqsbar_i;
  input [1:0] dm_i;
  input ri_i, ts_i, ck_i, cke_i, csbar_i, rasbar_i, casbar_i, webar_i, odt_i;
  output ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad,
         webar_pad, odt_pad;
  wire   SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24;

  SSTL18DDR2DIFF ck_sstl ( .PAD(ck_pad), .PADN(ckbar_pad), .Z(
        SYNOPSYS_UNCONNECTED_1), .A(ck_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_42 cke_sstl ( .PAD(cke_pad), .Z(SYNOPSYS_UNCONNECTED_2), .A(cke_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_41 casbar_sstl ( .PAD(casbar_pad), .Z(SYNOPSYS_UNCONNECTED_3), 
        .A(casbar_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_40 rasbar_sstl ( .PAD(rasbar_pad), .Z(SYNOPSYS_UNCONNECTED_4), 
        .A(rasbar_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_39 csbar_sstl ( .PAD(csbar_pad), .Z(SYNOPSYS_UNCONNECTED_5), .A(
        csbar_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_38 webar_sstl ( .PAD(webar_pad), .Z(SYNOPSYS_UNCONNECTED_6), .A(
        webar_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_37 odt_sstl ( .PAD(odt_pad), .Z(SYNOPSYS_UNCONNECTED_7), .A(odt_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_36 BA_0__sstl_ba ( .PAD(ba_pad[0]), .Z(SYNOPSYS_UNCONNECTED_8), 
        .A(ba_i[0]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_35 BA_1__sstl_ba ( .PAD(ba_pad[1]), .Z(SYNOPSYS_UNCONNECTED_9), 
        .A(ba_i[1]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_34 A_0__sstl_a ( .PAD(a_pad[0]), .Z(SYNOPSYS_UNCONNECTED_10), .A(
        a_i[0]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_33 A_1__sstl_a ( .PAD(a_pad[1]), .Z(SYNOPSYS_UNCONNECTED_11), .A(
        a_i[1]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_32 A_2__sstl_a ( .PAD(a_pad[2]), .Z(SYNOPSYS_UNCONNECTED_12), .A(
        a_i[2]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_31 A_3__sstl_a ( .PAD(a_pad[3]), .Z(SYNOPSYS_UNCONNECTED_13), .A(
        a_i[3]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_30 A_4__sstl_a ( .PAD(a_pad[4]), .Z(SYNOPSYS_UNCONNECTED_14), .A(
        a_i[4]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_29 A_5__sstl_a ( .PAD(a_pad[5]), .Z(SYNOPSYS_UNCONNECTED_15), .A(
        a_i[5]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_28 A_6__sstl_a ( .PAD(a_pad[6]), .Z(SYNOPSYS_UNCONNECTED_16), .A(
        a_i[6]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_27 A_7__sstl_a ( .PAD(a_pad[7]), .Z(SYNOPSYS_UNCONNECTED_17), .A(
        a_i[7]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_26 A_8__sstl_a ( .PAD(a_pad[8]), .Z(SYNOPSYS_UNCONNECTED_18), .A(
        a_i[8]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_25 A_9__sstl_a ( .PAD(a_pad[9]), .Z(SYNOPSYS_UNCONNECTED_19), .A(
        a_i[9]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_24 A_10__sstl_a ( .PAD(a_pad[10]), .Z(SYNOPSYS_UNCONNECTED_20), 
        .A(a_i[10]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_23 A_11__sstl_a ( .PAD(a_pad[11]), .Z(SYNOPSYS_UNCONNECTED_21), 
        .A(a_i[11]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_22 A_12__sstl_a ( .PAD(a_pad[12]), .Z(SYNOPSYS_UNCONNECTED_22), 
        .A(a_i[12]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_21 DQ_0__sstl_dq ( .PAD(dq_pad[0]), .Z(dq_o[0]), .A(dq_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_20 DQ_1__sstl_dq ( .PAD(dq_pad[1]), .Z(dq_o[1]), .A(dq_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_19 DQ_2__sstl_dq ( .PAD(dq_pad[2]), .Z(dq_o[2]), .A(dq_i[2]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_18 DQ_3__sstl_dq ( .PAD(dq_pad[3]), .Z(dq_o[3]), .A(dq_i[3]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_17 DQ_4__sstl_dq ( .PAD(dq_pad[4]), .Z(dq_o[4]), .A(dq_i[4]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_16 DQ_5__sstl_dq ( .PAD(dq_pad[5]), .Z(dq_o[5]), .A(dq_i[5]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_15 DQ_6__sstl_dq ( .PAD(dq_pad[6]), .Z(dq_o[6]), .A(dq_i[6]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_14 DQ_7__sstl_dq ( .PAD(dq_pad[7]), .Z(dq_o[7]), .A(dq_i[7]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_13 DQ_8__sstl_dq ( .PAD(dq_pad[8]), .Z(dq_o[8]), .A(dq_i[8]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_12 DQ_9__sstl_dq ( .PAD(dq_pad[9]), .Z(dq_o[9]), .A(dq_i[9]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_11 DQ_10__sstl_dq ( .PAD(dq_pad[10]), .Z(dq_o[10]), .A(dq_i[10]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_10 DQ_11__sstl_dq ( .PAD(dq_pad[11]), .Z(dq_o[11]), .A(dq_i[11]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_9 DQ_12__sstl_dq ( .PAD(dq_pad[12]), .Z(dq_o[12]), .A(dq_i[12]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_8 DQ_13__sstl_dq ( .PAD(dq_pad[13]), .Z(dq_o[13]), .A(dq_i[13]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_7 DQ_14__sstl_dq ( .PAD(dq_pad[14]), .Z(dq_o[14]), .A(dq_i[14]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_6 DQ_15__sstl_dq ( .PAD(dq_pad[15]), .Z(dq_o[15]), .A(dq_i[15]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_5 DQS_0__sstl_dqs ( .PAD(dqs_pad[0]), .Z(dqs_o[0]), .A(dqs_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_4 DQS_1__sstl_dqs ( .PAD(dqs_pad[1]), .Z(dqs_o[1]), .A(dqs_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_3 DQSBAR_0__sstl_dqsbar ( .PAD(dqsbar_pad[0]), .Z(dqsbar_o[0]), 
        .A(dqsbar_i[0]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_2 DQSBAR_1__sstl_dqsbar ( .PAD(dqsbar_pad[1]), .Z(dqsbar_o[1]), 
        .A(dqsbar_i[1]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR2_1 DM_0__sstl_dm ( .PAD(dm_pad[0]), .Z(SYNOPSYS_UNCONNECTED_23), 
        .A(dm_i[0]), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR2_0 DM_1__sstl_dm ( .PAD(dm_pad[1]), .Z(SYNOPSYS_UNCONNECTED_24), 
        .A(dm_i[1]), .RI(1'b0), .TS(1'b1) );
endmodule


module ddr2_init_engine ( ready, csbar, rasbar, casbar, webar, ba, a, odt, 
        ts_con, cke, clk, reset, init, ck );
  output [1:0] ba;
  output [12:0] a;
  input clk, reset, init, ck;
  output ready, csbar, rasbar, casbar, webar, odt, ts_con, cke;
  wire   flag, RESET, INIT, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n1, n2, n3, n4, n5, n6, n7, n8, n9, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45;
  wire   [16:0] counter;
  assign csbar = 1'b0;
  assign a[12] = 1'b0;
  assign a[11] = 1'b0;
  assign a[6] = 1'b0;
  assign ts_con = 1'b0;

  DFFPOSX1 RESET_reg ( .D(reset), .CLK(clk), .Q(RESET) );
  DFFPOSX1 INIT_reg ( .D(init), .CLK(clk), .Q(INIT) );
  DFFPOSX1 flag_reg ( .D(n659), .CLK(clk), .Q(flag) );
  DFFPOSX1 counter_reg_0_ ( .D(n658), .CLK(clk), .Q(counter[0]) );
  DFFPOSX1 counter_reg_1_ ( .D(n657), .CLK(clk), .Q(counter[1]) );
  DFFPOSX1 counter_reg_2_ ( .D(n656), .CLK(clk), .Q(counter[2]) );
  DFFPOSX1 counter_reg_3_ ( .D(n655), .CLK(clk), .Q(counter[3]) );
  DFFPOSX1 counter_reg_4_ ( .D(n654), .CLK(clk), .Q(counter[4]) );
  DFFPOSX1 counter_reg_5_ ( .D(n653), .CLK(clk), .Q(counter[5]) );
  DFFPOSX1 counter_reg_6_ ( .D(n652), .CLK(clk), .Q(counter[6]) );
  DFFPOSX1 counter_reg_7_ ( .D(n651), .CLK(clk), .Q(counter[7]) );
  DFFPOSX1 counter_reg_8_ ( .D(n650), .CLK(clk), .Q(counter[8]) );
  DFFPOSX1 counter_reg_9_ ( .D(n649), .CLK(clk), .Q(counter[9]) );
  DFFPOSX1 counter_reg_10_ ( .D(n648), .CLK(clk), .Q(counter[10]) );
  DFFPOSX1 counter_reg_11_ ( .D(n647), .CLK(clk), .Q(counter[11]) );
  DFFPOSX1 counter_reg_12_ ( .D(n646), .CLK(clk), .Q(counter[12]) );
  DFFPOSX1 counter_reg_13_ ( .D(n645), .CLK(clk), .Q(counter[13]) );
  DFFPOSX1 counter_reg_14_ ( .D(n644), .CLK(clk), .Q(counter[14]) );
  DFFPOSX1 counter_reg_15_ ( .D(n643), .CLK(clk), .Q(counter[15]) );
  DFFPOSX1 counter_reg_16_ ( .D(n642), .CLK(clk), .Q(counter[16]) );
  DFFPOSX1 ready_reg ( .D(n641), .CLK(clk), .Q(ready) );
  DFFPOSX1 casbar_reg ( .D(n640), .CLK(clk), .Q(casbar) );
  DFFPOSX1 webar_reg ( .D(n639), .CLK(clk), .Q(webar) );
  DFFPOSX1 rasbar_reg ( .D(n638), .CLK(clk), .Q(rasbar) );
  DFFPOSX1 cke_reg ( .D(n637), .CLK(clk), .Q(cke) );
  DFFPOSX1 odt_reg ( .D(n636), .CLK(clk), .Q(odt) );
  DFFPOSX1 a_reg_10_ ( .D(n635), .CLK(clk), .Q(a[10]) );
  DFFPOSX1 a_reg_9_ ( .D(n634), .CLK(clk), .Q(a[9]) );
  DFFPOSX1 a_reg_8_ ( .D(n633), .CLK(clk), .Q(a[8]) );
  DFFPOSX1 a_reg_7_ ( .D(n632), .CLK(clk), .Q(a[7]) );
  DFFPOSX1 a_reg_5_ ( .D(n631), .CLK(clk), .Q(a[5]) );
  DFFPOSX1 a_reg_4_ ( .D(n630), .CLK(clk), .Q(a[4]) );
  DFFPOSX1 a_reg_3_ ( .D(n629), .CLK(clk), .Q(a[3]) );
  DFFPOSX1 a_reg_2_ ( .D(n628), .CLK(clk), .Q(a[2]) );
  DFFPOSX1 a_reg_1_ ( .D(n627), .CLK(clk), .Q(a[1]) );
  DFFPOSX1 a_reg_0_ ( .D(n626), .CLK(clk), .Q(a[0]) );
  DFFPOSX1 ba_reg_1_ ( .D(n625), .CLK(clk), .Q(ba[1]) );
  DFFPOSX1 ba_reg_0_ ( .D(n624), .CLK(clk), .Q(ba[0]) );
  AOI21X1 U4 ( .A(ba[0]), .B(n453), .C(n454), .Y(n452) );
  OAI21X1 U5 ( .A(n455), .B(n456), .C(n457), .Y(n454) );
  OAI21X1 U6 ( .A(n458), .B(n456), .C(n459), .Y(n625) );
  NAND2X1 U7 ( .A(ba[1]), .B(n453), .Y(n459) );
  NAND3X1 U8 ( .A(n460), .B(n461), .C(n462), .Y(n456) );
  OAI21X1 U9 ( .A(n461), .B(n463), .C(n464), .Y(n626) );
  OAI21X1 U11 ( .A(n461), .B(n465), .C(n464), .Y(n627) );
  OAI21X1 U13 ( .A(n466), .B(n467), .C(n468), .Y(n628) );
  NAND2X1 U14 ( .A(a[2]), .B(n453), .Y(n468) );
  NAND2X1 U15 ( .A(n469), .B(n461), .Y(n467) );
  OAI21X1 U16 ( .A(n461), .B(n470), .C(n457), .Y(n629) );
  NAND2X1 U17 ( .A(n471), .B(n461), .Y(n457) );
  OAI21X1 U19 ( .A(n461), .B(n472), .C(n464), .Y(n630) );
  OAI21X1 U21 ( .A(n461), .B(n473), .C(n464), .Y(n631) );
  NAND3X1 U22 ( .A(n461), .B(n474), .C(n460), .Y(n464) );
  OAI21X1 U25 ( .A(n475), .B(n476), .C(n477), .Y(n632) );
  AOI21X1 U28 ( .A(a[8]), .B(n479), .C(n480), .Y(n478) );
  OAI21X1 U29 ( .A(n481), .B(n482), .C(n477), .Y(n480) );
  NAND2X1 U30 ( .A(n471), .B(n475), .Y(n477) );
  NAND2X1 U32 ( .A(n483), .B(n460), .Y(n466) );
  NAND2X1 U33 ( .A(n460), .B(n475), .Y(n482) );
  OAI21X1 U34 ( .A(n484), .B(n485), .C(n486), .Y(n634) );
  NAND2X1 U35 ( .A(a[9]), .B(n479), .Y(n486) );
  NAND2X1 U37 ( .A(n475), .B(n487), .Y(n485) );
  OAI21X1 U38 ( .A(n488), .B(n489), .C(n453), .Y(n475) );
  NAND2X1 U39 ( .A(n490), .B(n491), .Y(n489) );
  NAND2X1 U40 ( .A(n492), .B(n493), .Y(n488) );
  OAI21X1 U41 ( .A(n484), .B(n494), .C(n495), .Y(n635) );
  NAND2X1 U42 ( .A(a[10]), .B(n496), .Y(n495) );
  OAI21X1 U44 ( .A(n487), .B(n498), .C(n497), .Y(n494) );
  OAI21X1 U45 ( .A(n499), .B(n500), .C(n453), .Y(n497) );
  AOI21X1 U46 ( .A(n501), .B(n492), .C(RESET), .Y(n453) );
  OAI21X1 U48 ( .A(n503), .B(n504), .C(n505), .Y(n636) );
  NAND2X1 U49 ( .A(odt), .B(n45), .Y(n505) );
  NAND2X1 U50 ( .A(n507), .B(n508), .Y(n504) );
  OAI21X1 U51 ( .A(n509), .B(n510), .C(n511), .Y(n637) );
  NAND2X1 U52 ( .A(cke), .B(n45), .Y(n511) );
  NAND2X1 U53 ( .A(n512), .B(n507), .Y(n510) );
  NAND2X1 U54 ( .A(n492), .B(n513), .Y(n509) );
  OAI21X1 U55 ( .A(n484), .B(n514), .C(n515), .Y(n638) );
  NAND2X1 U56 ( .A(rasbar), .B(n516), .Y(n515) );
  NAND2X1 U57 ( .A(n517), .B(n518), .Y(n514) );
  OAI21X1 U58 ( .A(n484), .B(n519), .C(n520), .Y(n639) );
  NAND2X1 U59 ( .A(webar), .B(n516), .Y(n520) );
  NAND2X1 U61 ( .A(n517), .B(n521), .Y(n519) );
  NAND2X1 U62 ( .A(n45), .B(n522), .Y(n517) );
  OAI21X1 U63 ( .A(n523), .B(n524), .C(n525), .Y(n640) );
  OAI21X1 U64 ( .A(n498), .B(n518), .C(n523), .Y(n525) );
  OAI21X1 U68 ( .A(n527), .B(n528), .C(n492), .Y(n522) );
  NAND2X1 U70 ( .A(n529), .B(n526), .Y(n521) );
  NOR2X1 U71 ( .A(n530), .B(n531), .Y(n526) );
  OAI21X1 U72 ( .A(counter[2]), .B(n532), .C(n533), .Y(n531) );
  OAI21X1 U73 ( .A(n534), .B(n535), .C(n536), .Y(n533) );
  OAI21X1 U74 ( .A(n537), .B(n538), .C(n539), .Y(n535) );
  NAND3X1 U75 ( .A(n540), .B(n541), .C(counter[7]), .Y(n539) );
  NAND2X1 U76 ( .A(counter[3]), .B(n513), .Y(n538) );
  OAI21X1 U77 ( .A(n542), .B(n543), .C(n544), .Y(n534) );
  NAND2X1 U78 ( .A(n545), .B(n546), .Y(n543) );
  AOI22X1 U79 ( .A(n547), .B(counter[1]), .C(n548), .D(n549), .Y(n532) );
  OAI21X1 U80 ( .A(n542), .B(n550), .C(n551), .Y(n548) );
  NAND2X1 U81 ( .A(counter[6]), .B(n469), .Y(n550) );
  NOR2X1 U82 ( .A(n552), .B(n553), .Y(n547) );
  OAI21X1 U83 ( .A(n554), .B(n555), .C(n556), .Y(n530) );
  AOI22X1 U84 ( .A(n557), .B(n490), .C(n558), .D(n559), .Y(n556) );
  NOR2X1 U86 ( .A(n561), .B(n493), .Y(n557) );
  AOI22X1 U87 ( .A(n562), .B(n483), .C(n507), .D(n508), .Y(n561) );
  NOR2X1 U88 ( .A(n560), .B(n563), .Y(n507) );
  AOI21X1 U89 ( .A(n536), .B(n469), .C(n564), .Y(n554) );
  OAI21X1 U90 ( .A(n565), .B(n560), .C(n566), .Y(n564) );
  AOI22X1 U91 ( .A(n567), .B(n568), .C(n569), .D(n570), .Y(n529) );
  NAND3X1 U93 ( .A(counter[8]), .B(n563), .C(n512), .Y(n544) );
  NAND3X1 U95 ( .A(n571), .B(counter[5]), .C(n572), .Y(n537) );
  NOR2X1 U96 ( .A(n508), .B(n546), .Y(n572) );
  NOR2X1 U97 ( .A(n565), .B(n546), .Y(n568) );
  NOR2X1 U98 ( .A(n542), .B(n560), .Y(n567) );
  NAND2X1 U99 ( .A(counter[2]), .B(counter[1]), .Y(n560) );
  OAI22X1 U100 ( .A(n502), .B(n553), .C(n458), .D(n555), .Y(n501) );
  AOI22X1 U101 ( .A(n536), .B(n540), .C(n570), .D(n469), .Y(n458) );
  NAND2X1 U103 ( .A(counter[1]), .B(n573), .Y(n455) );
  AOI22X1 U105 ( .A(n474), .B(counter[1]), .C(n575), .D(n483), .Y(n502) );
  AOI22X1 U107 ( .A(n469), .B(counter[7]), .C(n576), .D(n562), .Y(n552) );
  NOR2X1 U108 ( .A(n563), .B(counter[4]), .Y(n469) );
  OAI21X1 U109 ( .A(n481), .B(n577), .C(n578), .Y(n474) );
  NAND3X1 U110 ( .A(n540), .B(n573), .C(counter[7]), .Y(n578) );
  NAND2X1 U111 ( .A(counter[2]), .B(n576), .Y(n577) );
  OAI21X1 U112 ( .A(n579), .B(n580), .C(n499), .Y(n527) );
  OAI21X1 U114 ( .A(n551), .B(n574), .C(n581), .Y(n498) );
  NAND3X1 U115 ( .A(n582), .B(n583), .C(n584), .Y(n581) );
  NOR2X1 U116 ( .A(counter[6]), .B(counter[2]), .Y(n584) );
  NAND3X1 U118 ( .A(counter[8]), .B(n493), .C(n571), .Y(n542) );
  NOR2X1 U119 ( .A(counter[9]), .B(counter[7]), .Y(n571) );
  NAND2X1 U120 ( .A(counter[2]), .B(n549), .Y(n574) );
  AOI21X1 U121 ( .A(n462), .B(n545), .C(n558), .Y(n551) );
  NAND3X1 U123 ( .A(n540), .B(counter[5]), .C(n490), .Y(n585) );
  NAND2X1 U125 ( .A(n563), .B(n508), .Y(n565) );
  NAND2X1 U127 ( .A(n541), .B(n576), .Y(n555) );
  NAND3X1 U129 ( .A(counter[8]), .B(counter[5]), .C(n586), .Y(n553) );
  NOR2X1 U130 ( .A(counter[9]), .B(counter[6]), .Y(n586) );
  NAND2X1 U131 ( .A(n491), .B(n493), .Y(n580) );
  NAND2X1 U133 ( .A(n583), .B(counter[2]), .Y(n566) );
  AND2X1 U134 ( .A(n545), .B(counter[1]), .Y(n583) );
  NOR2X1 U135 ( .A(n508), .B(n563), .Y(n545) );
  OAI21X1 U136 ( .A(n503), .B(n587), .C(n588), .Y(n641) );
  NAND2X1 U137 ( .A(ready), .B(n45), .Y(n588) );
  NAND2X1 U138 ( .A(n562), .B(n483), .Y(n587) );
  NOR2X1 U139 ( .A(counter[1]), .B(counter[2]), .Y(n483) );
  NAND2X1 U141 ( .A(counter[4]), .B(n563), .Y(n481) );
  NAND3X1 U142 ( .A(n492), .B(counter[5]), .C(n490), .Y(n503) );
  NAND3X1 U144 ( .A(counter[7]), .B(n513), .C(n589), .Y(n579) );
  NOR2X1 U145 ( .A(n546), .B(n590), .Y(n589) );
  NAND3X1 U147 ( .A(n591), .B(n592), .C(n593), .Y(n500) );
  NOR2X1 U148 ( .A(n594), .B(n595), .Y(n593) );
  NAND2X1 U149 ( .A(n460), .B(n596), .Y(n595) );
  NAND3X1 U151 ( .A(n597), .B(n598), .C(n599), .Y(n594) );
  NOR2X1 U152 ( .A(n600), .B(n601), .Y(n592) );
  NOR2X1 U153 ( .A(n602), .B(n603), .Y(n591) );
  INVX2 U3 ( .A(n452), .Y(n624) );
  INVX2 U10 ( .A(a[0]), .Y(n463) );
  INVX2 U12 ( .A(a[1]), .Y(n465) );
  INVX2 U18 ( .A(a[3]), .Y(n470) );
  INVX2 U20 ( .A(a[4]), .Y(n472) );
  INVX2 U23 ( .A(a[5]), .Y(n473) );
  INVX2 U26 ( .A(a[7]), .Y(n476) );
  INVX2 U27 ( .A(n478), .Y(n633) );
  INVX2 U31 ( .A(n466), .Y(n471) );
  INVX2 U36 ( .A(n475), .Y(n479) );
  INVX2 U43 ( .A(n497), .Y(n496) );
  INVX2 U47 ( .A(n502), .Y(n487) );
  INVX2 U60 ( .A(n517), .Y(n516) );
  INVX2 U65 ( .A(n526), .Y(n518) );
  INVX2 U66 ( .A(casbar), .Y(n524) );
  INVX2 U67 ( .A(n522), .Y(n523) );
  OR2X2 U69 ( .A(n501), .B(n521), .Y(n528) );
  INVX2 U85 ( .A(n560), .Y(n559) );
  INVX2 U92 ( .A(n544), .Y(n569) );
  INVX2 U94 ( .A(n537), .Y(n512) );
  INVX2 U102 ( .A(n455), .Y(n570) );
  INVX2 U104 ( .A(n574), .Y(n536) );
  INVX2 U106 ( .A(n552), .Y(n575) );
  INVX2 U113 ( .A(n498), .Y(n499) );
  INVX2 U117 ( .A(n542), .Y(n582) );
  INVX2 U122 ( .A(n585), .Y(n558) );
  INVX2 U124 ( .A(n565), .Y(n540) );
  INVX2 U126 ( .A(n555), .Y(n462) );
  INVX2 U128 ( .A(n553), .Y(n541) );
  INVX2 U132 ( .A(n566), .Y(n491) );
  INVX2 U140 ( .A(n481), .Y(n562) );
  INVX2 U143 ( .A(n579), .Y(n490) );
  INVX2 U146 ( .A(n500), .Y(n492) );
  INVX2 U150 ( .A(n484), .Y(n460) );
  INVX2 U174 ( .A(counter[10]), .Y(n600) );
  INVX2 U177 ( .A(counter[9]), .Y(n590) );
  INVX2 U180 ( .A(counter[8]), .Y(n513) );
  INVX2 U183 ( .A(counter[7]), .Y(n576) );
  INVX2 U186 ( .A(counter[6]), .Y(n546) );
  INVX2 U189 ( .A(counter[5]), .Y(n493) );
  INVX2 U192 ( .A(counter[4]), .Y(n508) );
  INVX2 U195 ( .A(counter[3]), .Y(n563) );
  INVX2 U198 ( .A(counter[2]), .Y(n573) );
  INVX2 U201 ( .A(counter[1]), .Y(n549) );
  INVX2 U205 ( .A(counter[0]), .Y(n596) );
  ddr2_init_engine_DW01_inc_1 add_103 ( .A(counter), .SUM({n26, n25, n24, n23, 
        n22, n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, n10}) );
  INVX2 U24 ( .A(n44), .Y(n38) );
  INVX2 U154 ( .A(n453), .Y(n461) );
  INVX2 U155 ( .A(RESET), .Y(n45) );
  NAND2X1 U156 ( .A(flag), .B(n45), .Y(n484) );
  INVX2 U157 ( .A(counter[13]), .Y(n602) );
  INVX2 U158 ( .A(counter[16]), .Y(n603) );
  INVX2 U159 ( .A(counter[11]), .Y(n601) );
  INVX2 U160 ( .A(counter[14]), .Y(n597) );
  INVX2 U161 ( .A(counter[15]), .Y(n598) );
  INVX2 U162 ( .A(counter[12]), .Y(n599) );
  INVX2 U163 ( .A(INIT), .Y(n1) );
  OAI21X1 U164 ( .A(RESET), .B(n1), .C(n484), .Y(n659) );
  INVX2 U165 ( .A(n659), .Y(n29) );
  NAND2X1 U166 ( .A(counter[16]), .B(n29), .Y(n3) );
  NAND2X1 U167 ( .A(flag), .B(n659), .Y(n44) );
  NAND2X1 U168 ( .A(n26), .B(n38), .Y(n2) );
  NAND2X1 U169 ( .A(n3), .B(n2), .Y(n642) );
  NAND2X1 U170 ( .A(counter[15]), .B(n29), .Y(n5) );
  NAND2X1 U171 ( .A(n25), .B(n38), .Y(n4) );
  NAND2X1 U172 ( .A(n5), .B(n4), .Y(n643) );
  NAND2X1 U173 ( .A(counter[14]), .B(n29), .Y(n7) );
  NAND2X1 U175 ( .A(n24), .B(n38), .Y(n6) );
  NAND2X1 U176 ( .A(n7), .B(n6), .Y(n644) );
  NAND2X1 U178 ( .A(counter[13]), .B(n29), .Y(n9) );
  NAND2X1 U179 ( .A(n23), .B(n38), .Y(n8) );
  NAND2X1 U181 ( .A(n9), .B(n8), .Y(n645) );
  NAND2X1 U182 ( .A(counter[12]), .B(n29), .Y(n28) );
  NAND2X1 U184 ( .A(n22), .B(n38), .Y(n27) );
  NAND2X1 U185 ( .A(n28), .B(n27), .Y(n646) );
  NAND2X1 U187 ( .A(counter[11]), .B(n29), .Y(n31) );
  NAND2X1 U188 ( .A(n21), .B(n38), .Y(n30) );
  NAND2X1 U190 ( .A(n31), .B(n30), .Y(n647) );
  NAND2X1 U191 ( .A(n20), .B(n38), .Y(n32) );
  OAI21X1 U193 ( .A(n659), .B(n600), .C(n32), .Y(n648) );
  NAND2X1 U194 ( .A(n19), .B(n38), .Y(n33) );
  OAI21X1 U196 ( .A(n659), .B(n590), .C(n33), .Y(n649) );
  NAND2X1 U197 ( .A(n18), .B(n38), .Y(n34) );
  OAI21X1 U199 ( .A(n659), .B(n513), .C(n34), .Y(n650) );
  NAND2X1 U200 ( .A(n17), .B(n38), .Y(n35) );
  OAI21X1 U202 ( .A(n659), .B(n576), .C(n35), .Y(n651) );
  NAND2X1 U203 ( .A(n16), .B(n38), .Y(n36) );
  OAI21X1 U204 ( .A(n659), .B(n546), .C(n36), .Y(n652) );
  NAND2X1 U206 ( .A(n15), .B(n38), .Y(n37) );
  OAI21X1 U207 ( .A(n659), .B(n493), .C(n37), .Y(n653) );
  NAND2X1 U208 ( .A(n14), .B(n38), .Y(n39) );
  OAI21X1 U209 ( .A(n659), .B(n508), .C(n39), .Y(n654) );
  INVX2 U210 ( .A(n13), .Y(n40) );
  OAI22X1 U216 ( .A(n659), .B(n563), .C(n44), .D(n40), .Y(n655) );
  INVX2 U217 ( .A(n12), .Y(n41) );
  OAI22X1 U218 ( .A(n659), .B(n573), .C(n44), .D(n41), .Y(n656) );
  INVX2 U219 ( .A(n11), .Y(n42) );
  OAI22X1 U220 ( .A(n659), .B(n549), .C(n44), .D(n42), .Y(n657) );
  INVX2 U221 ( .A(n10), .Y(n43) );
  OAI22X1 U222 ( .A(n659), .B(n596), .C(n44), .D(n43), .Y(n658) );
endmodule


module FIFO_DEPTH_P26_WIDTH41 ( clk, reset, data_in, put, get, data_out, empty, 
        full, fillcount );
  input [40:0] data_in;
  output [40:0] data_out;
  output [6:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   n13, n14, n15, n16, n17, n18, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7955, n7956, n7957, n7958, n7998, n7999, n8000, n8040,
         n8041, n8042, n8082, n8083, n8084, n8085, n8125, n8126, n8127, n8128,
         n8168, n8169, n8170, n8171, n8211, n8212, n8213, n8214, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10637, n10638, n10678, n10679, n10719, n10720, n10760,
         n10761, n10801, n10802, n10842, n10843, n10883, n10884, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556;
  wire   [5:0] wr_ptr;
  wire   [2623:0] arr;

  DFFPOSX1 fillcount_reg_0_ ( .D(n10938), .CLK(clk), .Q(fillcount[0]) );
  DFFPOSX1 fillcount_reg_1_ ( .D(n10937), .CLK(clk), .Q(fillcount[1]) );
  DFFPOSX1 fillcount_reg_6_ ( .D(n10936), .CLK(clk), .Q(fillcount[6]) );
  DFFPOSX1 fillcount_reg_2_ ( .D(n10935), .CLK(clk), .Q(fillcount[2]) );
  DFFPOSX1 fillcount_reg_3_ ( .D(n10934), .CLK(clk), .Q(fillcount[3]) );
  DFFPOSX1 fillcount_reg_4_ ( .D(n10933), .CLK(clk), .Q(fillcount[4]) );
  DFFPOSX1 fillcount_reg_5_ ( .D(n10932), .CLK(clk), .Q(fillcount[5]) );
  DFFPOSX1 wr_ptr_reg_0_ ( .D(n10931), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n10930), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n10929), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n10928), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n10927), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 wr_ptr_reg_5_ ( .D(n10926), .CLK(clk), .Q(wr_ptr[5]) );
  DFFPOSX1 arr_reg_63__40_ ( .D(n10925), .CLK(clk), .Q(arr[2623]) );
  DFFPOSX1 arr_reg_63__39_ ( .D(n10924), .CLK(clk), .Q(arr[2622]) );
  DFFPOSX1 arr_reg_63__38_ ( .D(n78), .CLK(clk), .Q(arr[2621]) );
  DFFPOSX1 arr_reg_63__37_ ( .D(n77), .CLK(clk), .Q(arr[2620]) );
  DFFPOSX1 arr_reg_63__36_ ( .D(n76), .CLK(clk), .Q(arr[2619]) );
  DFFPOSX1 arr_reg_63__35_ ( .D(n75), .CLK(clk), .Q(arr[2618]) );
  DFFPOSX1 arr_reg_63__34_ ( .D(n74), .CLK(clk), .Q(arr[2617]) );
  DFFPOSX1 arr_reg_63__33_ ( .D(n73), .CLK(clk), .Q(arr[2616]) );
  DFFPOSX1 arr_reg_63__32_ ( .D(n72), .CLK(clk), .Q(arr[2615]) );
  DFFPOSX1 arr_reg_63__31_ ( .D(n71), .CLK(clk), .Q(arr[2614]) );
  DFFPOSX1 arr_reg_63__30_ ( .D(n70), .CLK(clk), .Q(arr[2613]) );
  DFFPOSX1 arr_reg_63__29_ ( .D(n227), .CLK(clk), .Q(arr[2612]) );
  DFFPOSX1 arr_reg_63__28_ ( .D(n226), .CLK(clk), .Q(arr[2611]) );
  DFFPOSX1 arr_reg_63__27_ ( .D(n225), .CLK(clk), .Q(arr[2610]) );
  DFFPOSX1 arr_reg_63__26_ ( .D(n224), .CLK(clk), .Q(arr[2609]) );
  DFFPOSX1 arr_reg_63__25_ ( .D(n223), .CLK(clk), .Q(arr[2608]) );
  DFFPOSX1 arr_reg_63__24_ ( .D(n222), .CLK(clk), .Q(arr[2607]) );
  DFFPOSX1 arr_reg_63__23_ ( .D(n221), .CLK(clk), .Q(arr[2606]) );
  DFFPOSX1 arr_reg_63__22_ ( .D(n220), .CLK(clk), .Q(arr[2605]) );
  DFFPOSX1 arr_reg_63__21_ ( .D(n219), .CLK(clk), .Q(arr[2604]) );
  DFFPOSX1 arr_reg_63__20_ ( .D(n218), .CLK(clk), .Q(arr[2603]) );
  DFFPOSX1 arr_reg_63__19_ ( .D(n217), .CLK(clk), .Q(arr[2602]) );
  DFFPOSX1 arr_reg_63__18_ ( .D(n216), .CLK(clk), .Q(arr[2601]) );
  DFFPOSX1 arr_reg_63__17_ ( .D(n215), .CLK(clk), .Q(arr[2600]) );
  DFFPOSX1 arr_reg_63__16_ ( .D(n214), .CLK(clk), .Q(arr[2599]) );
  DFFPOSX1 arr_reg_63__15_ ( .D(n213), .CLK(clk), .Q(arr[2598]) );
  DFFPOSX1 arr_reg_63__14_ ( .D(n212), .CLK(clk), .Q(arr[2597]) );
  DFFPOSX1 arr_reg_63__13_ ( .D(n211), .CLK(clk), .Q(arr[2596]) );
  DFFPOSX1 arr_reg_63__12_ ( .D(n331), .CLK(clk), .Q(arr[2595]) );
  DFFPOSX1 arr_reg_63__11_ ( .D(n330), .CLK(clk), .Q(arr[2594]) );
  DFFPOSX1 arr_reg_63__10_ ( .D(n329), .CLK(clk), .Q(arr[2593]) );
  DFFPOSX1 arr_reg_63__9_ ( .D(n328), .CLK(clk), .Q(arr[2592]) );
  DFFPOSX1 arr_reg_63__8_ ( .D(n327), .CLK(clk), .Q(arr[2591]) );
  DFFPOSX1 arr_reg_63__7_ ( .D(n326), .CLK(clk), .Q(arr[2590]) );
  DFFPOSX1 arr_reg_63__6_ ( .D(n325), .CLK(clk), .Q(arr[2589]) );
  DFFPOSX1 arr_reg_63__5_ ( .D(n324), .CLK(clk), .Q(arr[2588]) );
  DFFPOSX1 arr_reg_63__4_ ( .D(n323), .CLK(clk), .Q(arr[2587]) );
  DFFPOSX1 arr_reg_63__3_ ( .D(n322), .CLK(clk), .Q(arr[2586]) );
  DFFPOSX1 arr_reg_63__2_ ( .D(n321), .CLK(clk), .Q(arr[2585]) );
  DFFPOSX1 arr_reg_63__1_ ( .D(n320), .CLK(clk), .Q(arr[2584]) );
  DFFPOSX1 arr_reg_63__0_ ( .D(n319), .CLK(clk), .Q(arr[2583]) );
  DFFPOSX1 arr_reg_62__40_ ( .D(n10884), .CLK(clk), .Q(arr[2582]) );
  DFFPOSX1 arr_reg_62__39_ ( .D(n10883), .CLK(clk), .Q(arr[2581]) );
  DFFPOSX1 arr_reg_62__38_ ( .D(n69), .CLK(clk), .Q(arr[2580]) );
  DFFPOSX1 arr_reg_62__37_ ( .D(n68), .CLK(clk), .Q(arr[2579]) );
  DFFPOSX1 arr_reg_62__36_ ( .D(n67), .CLK(clk), .Q(arr[2578]) );
  DFFPOSX1 arr_reg_62__35_ ( .D(n66), .CLK(clk), .Q(arr[2577]) );
  DFFPOSX1 arr_reg_62__34_ ( .D(n65), .CLK(clk), .Q(arr[2576]) );
  DFFPOSX1 arr_reg_62__33_ ( .D(n64), .CLK(clk), .Q(arr[2575]) );
  DFFPOSX1 arr_reg_62__32_ ( .D(n63), .CLK(clk), .Q(arr[2574]) );
  DFFPOSX1 arr_reg_62__31_ ( .D(n62), .CLK(clk), .Q(arr[2573]) );
  DFFPOSX1 arr_reg_62__30_ ( .D(n61), .CLK(clk), .Q(arr[2572]) );
  DFFPOSX1 arr_reg_62__29_ ( .D(n210), .CLK(clk), .Q(arr[2571]) );
  DFFPOSX1 arr_reg_62__28_ ( .D(n209), .CLK(clk), .Q(arr[2570]) );
  DFFPOSX1 arr_reg_62__27_ ( .D(n208), .CLK(clk), .Q(arr[2569]) );
  DFFPOSX1 arr_reg_62__26_ ( .D(n207), .CLK(clk), .Q(arr[2568]) );
  DFFPOSX1 arr_reg_62__25_ ( .D(n206), .CLK(clk), .Q(arr[2567]) );
  DFFPOSX1 arr_reg_62__24_ ( .D(n205), .CLK(clk), .Q(arr[2566]) );
  DFFPOSX1 arr_reg_62__23_ ( .D(n204), .CLK(clk), .Q(arr[2565]) );
  DFFPOSX1 arr_reg_62__22_ ( .D(n203), .CLK(clk), .Q(arr[2564]) );
  DFFPOSX1 arr_reg_62__21_ ( .D(n202), .CLK(clk), .Q(arr[2563]) );
  DFFPOSX1 arr_reg_62__20_ ( .D(n201), .CLK(clk), .Q(arr[2562]) );
  DFFPOSX1 arr_reg_62__19_ ( .D(n200), .CLK(clk), .Q(arr[2561]) );
  DFFPOSX1 arr_reg_62__18_ ( .D(n199), .CLK(clk), .Q(arr[2560]) );
  DFFPOSX1 arr_reg_62__17_ ( .D(n198), .CLK(clk), .Q(arr[2559]) );
  DFFPOSX1 arr_reg_62__16_ ( .D(n197), .CLK(clk), .Q(arr[2558]) );
  DFFPOSX1 arr_reg_62__15_ ( .D(n196), .CLK(clk), .Q(arr[2557]) );
  DFFPOSX1 arr_reg_62__14_ ( .D(n195), .CLK(clk), .Q(arr[2556]) );
  DFFPOSX1 arr_reg_62__13_ ( .D(n194), .CLK(clk), .Q(arr[2555]) );
  DFFPOSX1 arr_reg_62__12_ ( .D(n318), .CLK(clk), .Q(arr[2554]) );
  DFFPOSX1 arr_reg_62__11_ ( .D(n317), .CLK(clk), .Q(arr[2553]) );
  DFFPOSX1 arr_reg_62__10_ ( .D(n316), .CLK(clk), .Q(arr[2552]) );
  DFFPOSX1 arr_reg_62__9_ ( .D(n315), .CLK(clk), .Q(arr[2551]) );
  DFFPOSX1 arr_reg_62__8_ ( .D(n314), .CLK(clk), .Q(arr[2550]) );
  DFFPOSX1 arr_reg_62__7_ ( .D(n313), .CLK(clk), .Q(arr[2549]) );
  DFFPOSX1 arr_reg_62__6_ ( .D(n312), .CLK(clk), .Q(arr[2548]) );
  DFFPOSX1 arr_reg_62__5_ ( .D(n311), .CLK(clk), .Q(arr[2547]) );
  DFFPOSX1 arr_reg_62__4_ ( .D(n310), .CLK(clk), .Q(arr[2546]) );
  DFFPOSX1 arr_reg_62__3_ ( .D(n309), .CLK(clk), .Q(arr[2545]) );
  DFFPOSX1 arr_reg_62__2_ ( .D(n308), .CLK(clk), .Q(arr[2544]) );
  DFFPOSX1 arr_reg_62__1_ ( .D(n307), .CLK(clk), .Q(arr[2543]) );
  DFFPOSX1 arr_reg_62__0_ ( .D(n306), .CLK(clk), .Q(arr[2542]) );
  DFFPOSX1 arr_reg_61__40_ ( .D(n10843), .CLK(clk), .Q(arr[2541]) );
  DFFPOSX1 arr_reg_61__39_ ( .D(n10842), .CLK(clk), .Q(arr[2540]) );
  DFFPOSX1 arr_reg_61__38_ ( .D(n60), .CLK(clk), .Q(arr[2539]) );
  DFFPOSX1 arr_reg_61__37_ ( .D(n59), .CLK(clk), .Q(arr[2538]) );
  DFFPOSX1 arr_reg_61__36_ ( .D(n58), .CLK(clk), .Q(arr[2537]) );
  DFFPOSX1 arr_reg_61__35_ ( .D(n57), .CLK(clk), .Q(arr[2536]) );
  DFFPOSX1 arr_reg_61__34_ ( .D(n56), .CLK(clk), .Q(arr[2535]) );
  DFFPOSX1 arr_reg_61__33_ ( .D(n55), .CLK(clk), .Q(arr[2534]) );
  DFFPOSX1 arr_reg_61__32_ ( .D(n54), .CLK(clk), .Q(arr[2533]) );
  DFFPOSX1 arr_reg_61__31_ ( .D(n53), .CLK(clk), .Q(arr[2532]) );
  DFFPOSX1 arr_reg_61__30_ ( .D(n52), .CLK(clk), .Q(arr[2531]) );
  DFFPOSX1 arr_reg_61__29_ ( .D(n193), .CLK(clk), .Q(arr[2530]) );
  DFFPOSX1 arr_reg_61__28_ ( .D(n192), .CLK(clk), .Q(arr[2529]) );
  DFFPOSX1 arr_reg_61__27_ ( .D(n191), .CLK(clk), .Q(arr[2528]) );
  DFFPOSX1 arr_reg_61__26_ ( .D(n190), .CLK(clk), .Q(arr[2527]) );
  DFFPOSX1 arr_reg_61__25_ ( .D(n189), .CLK(clk), .Q(arr[2526]) );
  DFFPOSX1 arr_reg_61__24_ ( .D(n188), .CLK(clk), .Q(arr[2525]) );
  DFFPOSX1 arr_reg_61__23_ ( .D(n187), .CLK(clk), .Q(arr[2524]) );
  DFFPOSX1 arr_reg_61__22_ ( .D(n186), .CLK(clk), .Q(arr[2523]) );
  DFFPOSX1 arr_reg_61__21_ ( .D(n185), .CLK(clk), .Q(arr[2522]) );
  DFFPOSX1 arr_reg_61__20_ ( .D(n184), .CLK(clk), .Q(arr[2521]) );
  DFFPOSX1 arr_reg_61__19_ ( .D(n183), .CLK(clk), .Q(arr[2520]) );
  DFFPOSX1 arr_reg_61__18_ ( .D(n182), .CLK(clk), .Q(arr[2519]) );
  DFFPOSX1 arr_reg_61__17_ ( .D(n181), .CLK(clk), .Q(arr[2518]) );
  DFFPOSX1 arr_reg_61__16_ ( .D(n180), .CLK(clk), .Q(arr[2517]) );
  DFFPOSX1 arr_reg_61__15_ ( .D(n179), .CLK(clk), .Q(arr[2516]) );
  DFFPOSX1 arr_reg_61__14_ ( .D(n178), .CLK(clk), .Q(arr[2515]) );
  DFFPOSX1 arr_reg_61__13_ ( .D(n177), .CLK(clk), .Q(arr[2514]) );
  DFFPOSX1 arr_reg_61__12_ ( .D(n305), .CLK(clk), .Q(arr[2513]) );
  DFFPOSX1 arr_reg_61__11_ ( .D(n304), .CLK(clk), .Q(arr[2512]) );
  DFFPOSX1 arr_reg_61__10_ ( .D(n303), .CLK(clk), .Q(arr[2511]) );
  DFFPOSX1 arr_reg_61__9_ ( .D(n302), .CLK(clk), .Q(arr[2510]) );
  DFFPOSX1 arr_reg_61__8_ ( .D(n301), .CLK(clk), .Q(arr[2509]) );
  DFFPOSX1 arr_reg_61__7_ ( .D(n300), .CLK(clk), .Q(arr[2508]) );
  DFFPOSX1 arr_reg_61__6_ ( .D(n299), .CLK(clk), .Q(arr[2507]) );
  DFFPOSX1 arr_reg_61__5_ ( .D(n298), .CLK(clk), .Q(arr[2506]) );
  DFFPOSX1 arr_reg_61__4_ ( .D(n297), .CLK(clk), .Q(arr[2505]) );
  DFFPOSX1 arr_reg_61__3_ ( .D(n296), .CLK(clk), .Q(arr[2504]) );
  DFFPOSX1 arr_reg_61__2_ ( .D(n295), .CLK(clk), .Q(arr[2503]) );
  DFFPOSX1 arr_reg_61__1_ ( .D(n294), .CLK(clk), .Q(arr[2502]) );
  DFFPOSX1 arr_reg_61__0_ ( .D(n293), .CLK(clk), .Q(arr[2501]) );
  DFFPOSX1 arr_reg_60__40_ ( .D(n10802), .CLK(clk), .Q(arr[2500]) );
  DFFPOSX1 arr_reg_60__39_ ( .D(n10801), .CLK(clk), .Q(arr[2499]) );
  DFFPOSX1 arr_reg_60__38_ ( .D(n51), .CLK(clk), .Q(arr[2498]) );
  DFFPOSX1 arr_reg_60__37_ ( .D(n50), .CLK(clk), .Q(arr[2497]) );
  DFFPOSX1 arr_reg_60__36_ ( .D(n49), .CLK(clk), .Q(arr[2496]) );
  DFFPOSX1 arr_reg_60__35_ ( .D(n48), .CLK(clk), .Q(arr[2495]) );
  DFFPOSX1 arr_reg_60__34_ ( .D(n47), .CLK(clk), .Q(arr[2494]) );
  DFFPOSX1 arr_reg_60__33_ ( .D(n46), .CLK(clk), .Q(arr[2493]) );
  DFFPOSX1 arr_reg_60__32_ ( .D(n45), .CLK(clk), .Q(arr[2492]) );
  DFFPOSX1 arr_reg_60__31_ ( .D(n44), .CLK(clk), .Q(arr[2491]) );
  DFFPOSX1 arr_reg_60__30_ ( .D(n43), .CLK(clk), .Q(arr[2490]) );
  DFFPOSX1 arr_reg_60__29_ ( .D(n176), .CLK(clk), .Q(arr[2489]) );
  DFFPOSX1 arr_reg_60__28_ ( .D(n175), .CLK(clk), .Q(arr[2488]) );
  DFFPOSX1 arr_reg_60__27_ ( .D(n174), .CLK(clk), .Q(arr[2487]) );
  DFFPOSX1 arr_reg_60__26_ ( .D(n173), .CLK(clk), .Q(arr[2486]) );
  DFFPOSX1 arr_reg_60__25_ ( .D(n172), .CLK(clk), .Q(arr[2485]) );
  DFFPOSX1 arr_reg_60__24_ ( .D(n171), .CLK(clk), .Q(arr[2484]) );
  DFFPOSX1 arr_reg_60__23_ ( .D(n170), .CLK(clk), .Q(arr[2483]) );
  DFFPOSX1 arr_reg_60__22_ ( .D(n169), .CLK(clk), .Q(arr[2482]) );
  DFFPOSX1 arr_reg_60__21_ ( .D(n168), .CLK(clk), .Q(arr[2481]) );
  DFFPOSX1 arr_reg_60__20_ ( .D(n167), .CLK(clk), .Q(arr[2480]) );
  DFFPOSX1 arr_reg_60__19_ ( .D(n166), .CLK(clk), .Q(arr[2479]) );
  DFFPOSX1 arr_reg_60__18_ ( .D(n165), .CLK(clk), .Q(arr[2478]) );
  DFFPOSX1 arr_reg_60__17_ ( .D(n164), .CLK(clk), .Q(arr[2477]) );
  DFFPOSX1 arr_reg_60__16_ ( .D(n163), .CLK(clk), .Q(arr[2476]) );
  DFFPOSX1 arr_reg_60__15_ ( .D(n162), .CLK(clk), .Q(arr[2475]) );
  DFFPOSX1 arr_reg_60__14_ ( .D(n161), .CLK(clk), .Q(arr[2474]) );
  DFFPOSX1 arr_reg_60__13_ ( .D(n160), .CLK(clk), .Q(arr[2473]) );
  DFFPOSX1 arr_reg_60__12_ ( .D(n292), .CLK(clk), .Q(arr[2472]) );
  DFFPOSX1 arr_reg_60__11_ ( .D(n291), .CLK(clk), .Q(arr[2471]) );
  DFFPOSX1 arr_reg_60__10_ ( .D(n290), .CLK(clk), .Q(arr[2470]) );
  DFFPOSX1 arr_reg_60__9_ ( .D(n289), .CLK(clk), .Q(arr[2469]) );
  DFFPOSX1 arr_reg_60__8_ ( .D(n288), .CLK(clk), .Q(arr[2468]) );
  DFFPOSX1 arr_reg_60__7_ ( .D(n287), .CLK(clk), .Q(arr[2467]) );
  DFFPOSX1 arr_reg_60__6_ ( .D(n286), .CLK(clk), .Q(arr[2466]) );
  DFFPOSX1 arr_reg_60__5_ ( .D(n285), .CLK(clk), .Q(arr[2465]) );
  DFFPOSX1 arr_reg_60__4_ ( .D(n284), .CLK(clk), .Q(arr[2464]) );
  DFFPOSX1 arr_reg_60__3_ ( .D(n283), .CLK(clk), .Q(arr[2463]) );
  DFFPOSX1 arr_reg_60__2_ ( .D(n282), .CLK(clk), .Q(arr[2462]) );
  DFFPOSX1 arr_reg_60__1_ ( .D(n281), .CLK(clk), .Q(arr[2461]) );
  DFFPOSX1 arr_reg_60__0_ ( .D(n280), .CLK(clk), .Q(arr[2460]) );
  DFFPOSX1 arr_reg_59__40_ ( .D(n10761), .CLK(clk), .Q(arr[2459]) );
  DFFPOSX1 arr_reg_59__39_ ( .D(n10760), .CLK(clk), .Q(arr[2458]) );
  DFFPOSX1 arr_reg_59__38_ ( .D(n42), .CLK(clk), .Q(arr[2457]) );
  DFFPOSX1 arr_reg_59__37_ ( .D(n41), .CLK(clk), .Q(arr[2456]) );
  DFFPOSX1 arr_reg_59__36_ ( .D(n40), .CLK(clk), .Q(arr[2455]) );
  DFFPOSX1 arr_reg_59__35_ ( .D(n39), .CLK(clk), .Q(arr[2454]) );
  DFFPOSX1 arr_reg_59__34_ ( .D(n38), .CLK(clk), .Q(arr[2453]) );
  DFFPOSX1 arr_reg_59__33_ ( .D(n37), .CLK(clk), .Q(arr[2452]) );
  DFFPOSX1 arr_reg_59__32_ ( .D(n36), .CLK(clk), .Q(arr[2451]) );
  DFFPOSX1 arr_reg_59__31_ ( .D(n35), .CLK(clk), .Q(arr[2450]) );
  DFFPOSX1 arr_reg_59__30_ ( .D(n34), .CLK(clk), .Q(arr[2449]) );
  DFFPOSX1 arr_reg_59__29_ ( .D(n159), .CLK(clk), .Q(arr[2448]) );
  DFFPOSX1 arr_reg_59__28_ ( .D(n158), .CLK(clk), .Q(arr[2447]) );
  DFFPOSX1 arr_reg_59__27_ ( .D(n157), .CLK(clk), .Q(arr[2446]) );
  DFFPOSX1 arr_reg_59__26_ ( .D(n156), .CLK(clk), .Q(arr[2445]) );
  DFFPOSX1 arr_reg_59__25_ ( .D(n155), .CLK(clk), .Q(arr[2444]) );
  DFFPOSX1 arr_reg_59__24_ ( .D(n154), .CLK(clk), .Q(arr[2443]) );
  DFFPOSX1 arr_reg_59__23_ ( .D(n153), .CLK(clk), .Q(arr[2442]) );
  DFFPOSX1 arr_reg_59__22_ ( .D(n152), .CLK(clk), .Q(arr[2441]) );
  DFFPOSX1 arr_reg_59__21_ ( .D(n151), .CLK(clk), .Q(arr[2440]) );
  DFFPOSX1 arr_reg_59__20_ ( .D(n150), .CLK(clk), .Q(arr[2439]) );
  DFFPOSX1 arr_reg_59__19_ ( .D(n149), .CLK(clk), .Q(arr[2438]) );
  DFFPOSX1 arr_reg_59__18_ ( .D(n148), .CLK(clk), .Q(arr[2437]) );
  DFFPOSX1 arr_reg_59__17_ ( .D(n147), .CLK(clk), .Q(arr[2436]) );
  DFFPOSX1 arr_reg_59__16_ ( .D(n146), .CLK(clk), .Q(arr[2435]) );
  DFFPOSX1 arr_reg_59__15_ ( .D(n145), .CLK(clk), .Q(arr[2434]) );
  DFFPOSX1 arr_reg_59__14_ ( .D(n144), .CLK(clk), .Q(arr[2433]) );
  DFFPOSX1 arr_reg_59__13_ ( .D(n143), .CLK(clk), .Q(arr[2432]) );
  DFFPOSX1 arr_reg_59__12_ ( .D(n279), .CLK(clk), .Q(arr[2431]) );
  DFFPOSX1 arr_reg_59__11_ ( .D(n278), .CLK(clk), .Q(arr[2430]) );
  DFFPOSX1 arr_reg_59__10_ ( .D(n277), .CLK(clk), .Q(arr[2429]) );
  DFFPOSX1 arr_reg_59__9_ ( .D(n276), .CLK(clk), .Q(arr[2428]) );
  DFFPOSX1 arr_reg_59__8_ ( .D(n275), .CLK(clk), .Q(arr[2427]) );
  DFFPOSX1 arr_reg_59__7_ ( .D(n274), .CLK(clk), .Q(arr[2426]) );
  DFFPOSX1 arr_reg_59__6_ ( .D(n273), .CLK(clk), .Q(arr[2425]) );
  DFFPOSX1 arr_reg_59__5_ ( .D(n272), .CLK(clk), .Q(arr[2424]) );
  DFFPOSX1 arr_reg_59__4_ ( .D(n271), .CLK(clk), .Q(arr[2423]) );
  DFFPOSX1 arr_reg_59__3_ ( .D(n270), .CLK(clk), .Q(arr[2422]) );
  DFFPOSX1 arr_reg_59__2_ ( .D(n269), .CLK(clk), .Q(arr[2421]) );
  DFFPOSX1 arr_reg_59__1_ ( .D(n268), .CLK(clk), .Q(arr[2420]) );
  DFFPOSX1 arr_reg_59__0_ ( .D(n267), .CLK(clk), .Q(arr[2419]) );
  DFFPOSX1 arr_reg_58__40_ ( .D(n10720), .CLK(clk), .Q(arr[2418]) );
  DFFPOSX1 arr_reg_58__39_ ( .D(n10719), .CLK(clk), .Q(arr[2417]) );
  DFFPOSX1 arr_reg_58__38_ ( .D(n33), .CLK(clk), .Q(arr[2416]) );
  DFFPOSX1 arr_reg_58__37_ ( .D(n32), .CLK(clk), .Q(arr[2415]) );
  DFFPOSX1 arr_reg_58__36_ ( .D(n31), .CLK(clk), .Q(arr[2414]) );
  DFFPOSX1 arr_reg_58__35_ ( .D(n30), .CLK(clk), .Q(arr[2413]) );
  DFFPOSX1 arr_reg_58__34_ ( .D(n29), .CLK(clk), .Q(arr[2412]) );
  DFFPOSX1 arr_reg_58__33_ ( .D(n28), .CLK(clk), .Q(arr[2411]) );
  DFFPOSX1 arr_reg_58__32_ ( .D(n27), .CLK(clk), .Q(arr[2410]) );
  DFFPOSX1 arr_reg_58__31_ ( .D(n26), .CLK(clk), .Q(arr[2409]) );
  DFFPOSX1 arr_reg_58__30_ ( .D(n25), .CLK(clk), .Q(arr[2408]) );
  DFFPOSX1 arr_reg_58__29_ ( .D(n142), .CLK(clk), .Q(arr[2407]) );
  DFFPOSX1 arr_reg_58__28_ ( .D(n141), .CLK(clk), .Q(arr[2406]) );
  DFFPOSX1 arr_reg_58__27_ ( .D(n140), .CLK(clk), .Q(arr[2405]) );
  DFFPOSX1 arr_reg_58__26_ ( .D(n139), .CLK(clk), .Q(arr[2404]) );
  DFFPOSX1 arr_reg_58__25_ ( .D(n138), .CLK(clk), .Q(arr[2403]) );
  DFFPOSX1 arr_reg_58__24_ ( .D(n137), .CLK(clk), .Q(arr[2402]) );
  DFFPOSX1 arr_reg_58__23_ ( .D(n136), .CLK(clk), .Q(arr[2401]) );
  DFFPOSX1 arr_reg_58__22_ ( .D(n135), .CLK(clk), .Q(arr[2400]) );
  DFFPOSX1 arr_reg_58__21_ ( .D(n134), .CLK(clk), .Q(arr[2399]) );
  DFFPOSX1 arr_reg_58__20_ ( .D(n133), .CLK(clk), .Q(arr[2398]) );
  DFFPOSX1 arr_reg_58__19_ ( .D(n132), .CLK(clk), .Q(arr[2397]) );
  DFFPOSX1 arr_reg_58__18_ ( .D(n131), .CLK(clk), .Q(arr[2396]) );
  DFFPOSX1 arr_reg_58__17_ ( .D(n130), .CLK(clk), .Q(arr[2395]) );
  DFFPOSX1 arr_reg_58__16_ ( .D(n129), .CLK(clk), .Q(arr[2394]) );
  DFFPOSX1 arr_reg_58__15_ ( .D(n128), .CLK(clk), .Q(arr[2393]) );
  DFFPOSX1 arr_reg_58__14_ ( .D(n127), .CLK(clk), .Q(arr[2392]) );
  DFFPOSX1 arr_reg_58__13_ ( .D(n126), .CLK(clk), .Q(arr[2391]) );
  DFFPOSX1 arr_reg_58__12_ ( .D(n266), .CLK(clk), .Q(arr[2390]) );
  DFFPOSX1 arr_reg_58__11_ ( .D(n265), .CLK(clk), .Q(arr[2389]) );
  DFFPOSX1 arr_reg_58__10_ ( .D(n264), .CLK(clk), .Q(arr[2388]) );
  DFFPOSX1 arr_reg_58__9_ ( .D(n263), .CLK(clk), .Q(arr[2387]) );
  DFFPOSX1 arr_reg_58__8_ ( .D(n262), .CLK(clk), .Q(arr[2386]) );
  DFFPOSX1 arr_reg_58__7_ ( .D(n261), .CLK(clk), .Q(arr[2385]) );
  DFFPOSX1 arr_reg_58__6_ ( .D(n260), .CLK(clk), .Q(arr[2384]) );
  DFFPOSX1 arr_reg_58__5_ ( .D(n259), .CLK(clk), .Q(arr[2383]) );
  DFFPOSX1 arr_reg_58__4_ ( .D(n258), .CLK(clk), .Q(arr[2382]) );
  DFFPOSX1 arr_reg_58__3_ ( .D(n257), .CLK(clk), .Q(arr[2381]) );
  DFFPOSX1 arr_reg_58__2_ ( .D(n256), .CLK(clk), .Q(arr[2380]) );
  DFFPOSX1 arr_reg_58__1_ ( .D(n255), .CLK(clk), .Q(arr[2379]) );
  DFFPOSX1 arr_reg_58__0_ ( .D(n254), .CLK(clk), .Q(arr[2378]) );
  DFFPOSX1 arr_reg_57__40_ ( .D(n10679), .CLK(clk), .Q(arr[2377]) );
  DFFPOSX1 arr_reg_57__39_ ( .D(n10678), .CLK(clk), .Q(arr[2376]) );
  DFFPOSX1 arr_reg_57__38_ ( .D(n24), .CLK(clk), .Q(arr[2375]) );
  DFFPOSX1 arr_reg_57__37_ ( .D(n23), .CLK(clk), .Q(arr[2374]) );
  DFFPOSX1 arr_reg_57__36_ ( .D(n22), .CLK(clk), .Q(arr[2373]) );
  DFFPOSX1 arr_reg_57__35_ ( .D(n21), .CLK(clk), .Q(arr[2372]) );
  DFFPOSX1 arr_reg_57__34_ ( .D(n20), .CLK(clk), .Q(arr[2371]) );
  DFFPOSX1 arr_reg_57__33_ ( .D(n19), .CLK(clk), .Q(arr[2370]) );
  DFFPOSX1 arr_reg_57__32_ ( .D(n12), .CLK(clk), .Q(arr[2369]) );
  DFFPOSX1 arr_reg_57__31_ ( .D(n11), .CLK(clk), .Q(arr[2368]) );
  DFFPOSX1 arr_reg_57__30_ ( .D(n10), .CLK(clk), .Q(arr[2367]) );
  DFFPOSX1 arr_reg_57__29_ ( .D(n125), .CLK(clk), .Q(arr[2366]) );
  DFFPOSX1 arr_reg_57__28_ ( .D(n124), .CLK(clk), .Q(arr[2365]) );
  DFFPOSX1 arr_reg_57__27_ ( .D(n123), .CLK(clk), .Q(arr[2364]) );
  DFFPOSX1 arr_reg_57__26_ ( .D(n122), .CLK(clk), .Q(arr[2363]) );
  DFFPOSX1 arr_reg_57__25_ ( .D(n121), .CLK(clk), .Q(arr[2362]) );
  DFFPOSX1 arr_reg_57__24_ ( .D(n120), .CLK(clk), .Q(arr[2361]) );
  DFFPOSX1 arr_reg_57__23_ ( .D(n119), .CLK(clk), .Q(arr[2360]) );
  DFFPOSX1 arr_reg_57__22_ ( .D(n118), .CLK(clk), .Q(arr[2359]) );
  DFFPOSX1 arr_reg_57__21_ ( .D(n117), .CLK(clk), .Q(arr[2358]) );
  DFFPOSX1 arr_reg_57__20_ ( .D(n116), .CLK(clk), .Q(arr[2357]) );
  DFFPOSX1 arr_reg_57__19_ ( .D(n115), .CLK(clk), .Q(arr[2356]) );
  DFFPOSX1 arr_reg_57__18_ ( .D(n114), .CLK(clk), .Q(arr[2355]) );
  DFFPOSX1 arr_reg_57__17_ ( .D(n113), .CLK(clk), .Q(arr[2354]) );
  DFFPOSX1 arr_reg_57__16_ ( .D(n112), .CLK(clk), .Q(arr[2353]) );
  DFFPOSX1 arr_reg_57__15_ ( .D(n111), .CLK(clk), .Q(arr[2352]) );
  DFFPOSX1 arr_reg_57__14_ ( .D(n110), .CLK(clk), .Q(arr[2351]) );
  DFFPOSX1 arr_reg_57__13_ ( .D(n109), .CLK(clk), .Q(arr[2350]) );
  DFFPOSX1 arr_reg_57__12_ ( .D(n253), .CLK(clk), .Q(arr[2349]) );
  DFFPOSX1 arr_reg_57__11_ ( .D(n252), .CLK(clk), .Q(arr[2348]) );
  DFFPOSX1 arr_reg_57__10_ ( .D(n251), .CLK(clk), .Q(arr[2347]) );
  DFFPOSX1 arr_reg_57__9_ ( .D(n250), .CLK(clk), .Q(arr[2346]) );
  DFFPOSX1 arr_reg_57__8_ ( .D(n249), .CLK(clk), .Q(arr[2345]) );
  DFFPOSX1 arr_reg_57__7_ ( .D(n248), .CLK(clk), .Q(arr[2344]) );
  DFFPOSX1 arr_reg_57__6_ ( .D(n247), .CLK(clk), .Q(arr[2343]) );
  DFFPOSX1 arr_reg_57__5_ ( .D(n246), .CLK(clk), .Q(arr[2342]) );
  DFFPOSX1 arr_reg_57__4_ ( .D(n245), .CLK(clk), .Q(arr[2341]) );
  DFFPOSX1 arr_reg_57__3_ ( .D(n244), .CLK(clk), .Q(arr[2340]) );
  DFFPOSX1 arr_reg_57__2_ ( .D(n243), .CLK(clk), .Q(arr[2339]) );
  DFFPOSX1 arr_reg_57__1_ ( .D(n242), .CLK(clk), .Q(arr[2338]) );
  DFFPOSX1 arr_reg_57__0_ ( .D(n241), .CLK(clk), .Q(arr[2337]) );
  DFFPOSX1 arr_reg_56__40_ ( .D(n10638), .CLK(clk), .Q(arr[2336]) );
  DFFPOSX1 arr_reg_56__39_ ( .D(n10637), .CLK(clk), .Q(arr[2335]) );
  DFFPOSX1 arr_reg_56__38_ ( .D(n9), .CLK(clk), .Q(arr[2334]) );
  DFFPOSX1 arr_reg_56__37_ ( .D(n8), .CLK(clk), .Q(arr[2333]) );
  DFFPOSX1 arr_reg_56__36_ ( .D(n7), .CLK(clk), .Q(arr[2332]) );
  DFFPOSX1 arr_reg_56__35_ ( .D(n6), .CLK(clk), .Q(arr[2331]) );
  DFFPOSX1 arr_reg_56__34_ ( .D(n5), .CLK(clk), .Q(arr[2330]) );
  DFFPOSX1 arr_reg_56__33_ ( .D(n4), .CLK(clk), .Q(arr[2329]) );
  DFFPOSX1 arr_reg_56__32_ ( .D(n3), .CLK(clk), .Q(arr[2328]) );
  DFFPOSX1 arr_reg_56__31_ ( .D(n2), .CLK(clk), .Q(arr[2327]) );
  DFFPOSX1 arr_reg_56__30_ ( .D(n1), .CLK(clk), .Q(arr[2326]) );
  DFFPOSX1 arr_reg_56__29_ ( .D(n108), .CLK(clk), .Q(arr[2325]) );
  DFFPOSX1 arr_reg_56__28_ ( .D(n107), .CLK(clk), .Q(arr[2324]) );
  DFFPOSX1 arr_reg_56__27_ ( .D(n106), .CLK(clk), .Q(arr[2323]) );
  DFFPOSX1 arr_reg_56__26_ ( .D(n105), .CLK(clk), .Q(arr[2322]) );
  DFFPOSX1 arr_reg_56__25_ ( .D(n104), .CLK(clk), .Q(arr[2321]) );
  DFFPOSX1 arr_reg_56__24_ ( .D(n103), .CLK(clk), .Q(arr[2320]) );
  DFFPOSX1 arr_reg_56__23_ ( .D(n102), .CLK(clk), .Q(arr[2319]) );
  DFFPOSX1 arr_reg_56__22_ ( .D(n101), .CLK(clk), .Q(arr[2318]) );
  DFFPOSX1 arr_reg_56__21_ ( .D(n100), .CLK(clk), .Q(arr[2317]) );
  DFFPOSX1 arr_reg_56__20_ ( .D(n99), .CLK(clk), .Q(arr[2316]) );
  DFFPOSX1 arr_reg_56__19_ ( .D(n85), .CLK(clk), .Q(arr[2315]) );
  DFFPOSX1 arr_reg_56__18_ ( .D(n84), .CLK(clk), .Q(arr[2314]) );
  DFFPOSX1 arr_reg_56__17_ ( .D(n83), .CLK(clk), .Q(arr[2313]) );
  DFFPOSX1 arr_reg_56__16_ ( .D(n82), .CLK(clk), .Q(arr[2312]) );
  DFFPOSX1 arr_reg_56__15_ ( .D(n81), .CLK(clk), .Q(arr[2311]) );
  DFFPOSX1 arr_reg_56__14_ ( .D(n80), .CLK(clk), .Q(arr[2310]) );
  DFFPOSX1 arr_reg_56__13_ ( .D(n79), .CLK(clk), .Q(arr[2309]) );
  DFFPOSX1 arr_reg_56__12_ ( .D(n240), .CLK(clk), .Q(arr[2308]) );
  DFFPOSX1 arr_reg_56__11_ ( .D(n239), .CLK(clk), .Q(arr[2307]) );
  DFFPOSX1 arr_reg_56__10_ ( .D(n238), .CLK(clk), .Q(arr[2306]) );
  DFFPOSX1 arr_reg_56__9_ ( .D(n237), .CLK(clk), .Q(arr[2305]) );
  DFFPOSX1 arr_reg_56__8_ ( .D(n236), .CLK(clk), .Q(arr[2304]) );
  DFFPOSX1 arr_reg_56__7_ ( .D(n235), .CLK(clk), .Q(arr[2303]) );
  DFFPOSX1 arr_reg_56__6_ ( .D(n234), .CLK(clk), .Q(arr[2302]) );
  DFFPOSX1 arr_reg_56__5_ ( .D(n233), .CLK(clk), .Q(arr[2301]) );
  DFFPOSX1 arr_reg_56__4_ ( .D(n232), .CLK(clk), .Q(arr[2300]) );
  DFFPOSX1 arr_reg_56__3_ ( .D(n231), .CLK(clk), .Q(arr[2299]) );
  DFFPOSX1 arr_reg_56__2_ ( .D(n230), .CLK(clk), .Q(arr[2298]) );
  DFFPOSX1 arr_reg_56__1_ ( .D(n229), .CLK(clk), .Q(arr[2297]) );
  DFFPOSX1 arr_reg_56__0_ ( .D(n228), .CLK(clk), .Q(arr[2296]) );
  DFFPOSX1 arr_reg_55__40_ ( .D(n10597), .CLK(clk), .Q(arr[2295]) );
  DFFPOSX1 arr_reg_55__39_ ( .D(n10596), .CLK(clk), .Q(arr[2294]) );
  DFFPOSX1 arr_reg_55__38_ ( .D(n10595), .CLK(clk), .Q(arr[2293]) );
  DFFPOSX1 arr_reg_55__37_ ( .D(n10594), .CLK(clk), .Q(arr[2292]) );
  DFFPOSX1 arr_reg_55__36_ ( .D(n10593), .CLK(clk), .Q(arr[2291]) );
  DFFPOSX1 arr_reg_55__35_ ( .D(n10592), .CLK(clk), .Q(arr[2290]) );
  DFFPOSX1 arr_reg_55__34_ ( .D(n10591), .CLK(clk), .Q(arr[2289]) );
  DFFPOSX1 arr_reg_55__33_ ( .D(n10590), .CLK(clk), .Q(arr[2288]) );
  DFFPOSX1 arr_reg_55__32_ ( .D(n10589), .CLK(clk), .Q(arr[2287]) );
  DFFPOSX1 arr_reg_55__31_ ( .D(n10588), .CLK(clk), .Q(arr[2286]) );
  DFFPOSX1 arr_reg_55__30_ ( .D(n10587), .CLK(clk), .Q(arr[2285]) );
  DFFPOSX1 arr_reg_55__29_ ( .D(n10586), .CLK(clk), .Q(arr[2284]) );
  DFFPOSX1 arr_reg_55__28_ ( .D(n10585), .CLK(clk), .Q(arr[2283]) );
  DFFPOSX1 arr_reg_55__27_ ( .D(n10584), .CLK(clk), .Q(arr[2282]) );
  DFFPOSX1 arr_reg_55__26_ ( .D(n10583), .CLK(clk), .Q(arr[2281]) );
  DFFPOSX1 arr_reg_55__25_ ( .D(n10582), .CLK(clk), .Q(arr[2280]) );
  DFFPOSX1 arr_reg_55__24_ ( .D(n10581), .CLK(clk), .Q(arr[2279]) );
  DFFPOSX1 arr_reg_55__23_ ( .D(n10580), .CLK(clk), .Q(arr[2278]) );
  DFFPOSX1 arr_reg_55__22_ ( .D(n10579), .CLK(clk), .Q(arr[2277]) );
  DFFPOSX1 arr_reg_55__21_ ( .D(n10578), .CLK(clk), .Q(arr[2276]) );
  DFFPOSX1 arr_reg_55__20_ ( .D(n10577), .CLK(clk), .Q(arr[2275]) );
  DFFPOSX1 arr_reg_55__19_ ( .D(n10576), .CLK(clk), .Q(arr[2274]) );
  DFFPOSX1 arr_reg_55__18_ ( .D(n10575), .CLK(clk), .Q(arr[2273]) );
  DFFPOSX1 arr_reg_55__17_ ( .D(n10574), .CLK(clk), .Q(arr[2272]) );
  DFFPOSX1 arr_reg_55__16_ ( .D(n10573), .CLK(clk), .Q(arr[2271]) );
  DFFPOSX1 arr_reg_55__15_ ( .D(n10572), .CLK(clk), .Q(arr[2270]) );
  DFFPOSX1 arr_reg_55__14_ ( .D(n10571), .CLK(clk), .Q(arr[2269]) );
  DFFPOSX1 arr_reg_55__13_ ( .D(n10570), .CLK(clk), .Q(arr[2268]) );
  DFFPOSX1 arr_reg_55__12_ ( .D(n10569), .CLK(clk), .Q(arr[2267]) );
  DFFPOSX1 arr_reg_55__11_ ( .D(n10568), .CLK(clk), .Q(arr[2266]) );
  DFFPOSX1 arr_reg_55__10_ ( .D(n10567), .CLK(clk), .Q(arr[2265]) );
  DFFPOSX1 arr_reg_55__9_ ( .D(n10566), .CLK(clk), .Q(arr[2264]) );
  DFFPOSX1 arr_reg_55__8_ ( .D(n10565), .CLK(clk), .Q(arr[2263]) );
  DFFPOSX1 arr_reg_55__7_ ( .D(n10564), .CLK(clk), .Q(arr[2262]) );
  DFFPOSX1 arr_reg_55__6_ ( .D(n10563), .CLK(clk), .Q(arr[2261]) );
  DFFPOSX1 arr_reg_55__5_ ( .D(n10562), .CLK(clk), .Q(arr[2260]) );
  DFFPOSX1 arr_reg_55__4_ ( .D(n10561), .CLK(clk), .Q(arr[2259]) );
  DFFPOSX1 arr_reg_55__3_ ( .D(n10560), .CLK(clk), .Q(arr[2258]) );
  DFFPOSX1 arr_reg_55__2_ ( .D(n10559), .CLK(clk), .Q(arr[2257]) );
  DFFPOSX1 arr_reg_55__1_ ( .D(n10558), .CLK(clk), .Q(arr[2256]) );
  DFFPOSX1 arr_reg_55__0_ ( .D(n10557), .CLK(clk), .Q(arr[2255]) );
  DFFPOSX1 arr_reg_54__40_ ( .D(n10556), .CLK(clk), .Q(arr[2254]) );
  DFFPOSX1 arr_reg_54__39_ ( .D(n10555), .CLK(clk), .Q(arr[2253]) );
  DFFPOSX1 arr_reg_54__38_ ( .D(n10554), .CLK(clk), .Q(arr[2252]) );
  DFFPOSX1 arr_reg_54__37_ ( .D(n10553), .CLK(clk), .Q(arr[2251]) );
  DFFPOSX1 arr_reg_54__36_ ( .D(n10552), .CLK(clk), .Q(arr[2250]) );
  DFFPOSX1 arr_reg_54__35_ ( .D(n10551), .CLK(clk), .Q(arr[2249]) );
  DFFPOSX1 arr_reg_54__34_ ( .D(n10550), .CLK(clk), .Q(arr[2248]) );
  DFFPOSX1 arr_reg_54__33_ ( .D(n10549), .CLK(clk), .Q(arr[2247]) );
  DFFPOSX1 arr_reg_54__32_ ( .D(n10548), .CLK(clk), .Q(arr[2246]) );
  DFFPOSX1 arr_reg_54__31_ ( .D(n10547), .CLK(clk), .Q(arr[2245]) );
  DFFPOSX1 arr_reg_54__30_ ( .D(n10546), .CLK(clk), .Q(arr[2244]) );
  DFFPOSX1 arr_reg_54__29_ ( .D(n10545), .CLK(clk), .Q(arr[2243]) );
  DFFPOSX1 arr_reg_54__28_ ( .D(n10544), .CLK(clk), .Q(arr[2242]) );
  DFFPOSX1 arr_reg_54__27_ ( .D(n10543), .CLK(clk), .Q(arr[2241]) );
  DFFPOSX1 arr_reg_54__26_ ( .D(n10542), .CLK(clk), .Q(arr[2240]) );
  DFFPOSX1 arr_reg_54__25_ ( .D(n10541), .CLK(clk), .Q(arr[2239]) );
  DFFPOSX1 arr_reg_54__24_ ( .D(n10540), .CLK(clk), .Q(arr[2238]) );
  DFFPOSX1 arr_reg_54__23_ ( .D(n10539), .CLK(clk), .Q(arr[2237]) );
  DFFPOSX1 arr_reg_54__22_ ( .D(n10538), .CLK(clk), .Q(arr[2236]) );
  DFFPOSX1 arr_reg_54__21_ ( .D(n10537), .CLK(clk), .Q(arr[2235]) );
  DFFPOSX1 arr_reg_54__20_ ( .D(n10536), .CLK(clk), .Q(arr[2234]) );
  DFFPOSX1 arr_reg_54__19_ ( .D(n10535), .CLK(clk), .Q(arr[2233]) );
  DFFPOSX1 arr_reg_54__18_ ( .D(n10534), .CLK(clk), .Q(arr[2232]) );
  DFFPOSX1 arr_reg_54__17_ ( .D(n10533), .CLK(clk), .Q(arr[2231]) );
  DFFPOSX1 arr_reg_54__16_ ( .D(n10532), .CLK(clk), .Q(arr[2230]) );
  DFFPOSX1 arr_reg_54__15_ ( .D(n10531), .CLK(clk), .Q(arr[2229]) );
  DFFPOSX1 arr_reg_54__14_ ( .D(n10530), .CLK(clk), .Q(arr[2228]) );
  DFFPOSX1 arr_reg_54__13_ ( .D(n10529), .CLK(clk), .Q(arr[2227]) );
  DFFPOSX1 arr_reg_54__12_ ( .D(n10528), .CLK(clk), .Q(arr[2226]) );
  DFFPOSX1 arr_reg_54__11_ ( .D(n10527), .CLK(clk), .Q(arr[2225]) );
  DFFPOSX1 arr_reg_54__10_ ( .D(n10526), .CLK(clk), .Q(arr[2224]) );
  DFFPOSX1 arr_reg_54__9_ ( .D(n10525), .CLK(clk), .Q(arr[2223]) );
  DFFPOSX1 arr_reg_54__8_ ( .D(n10524), .CLK(clk), .Q(arr[2222]) );
  DFFPOSX1 arr_reg_54__7_ ( .D(n10523), .CLK(clk), .Q(arr[2221]) );
  DFFPOSX1 arr_reg_54__6_ ( .D(n10522), .CLK(clk), .Q(arr[2220]) );
  DFFPOSX1 arr_reg_54__5_ ( .D(n10521), .CLK(clk), .Q(arr[2219]) );
  DFFPOSX1 arr_reg_54__4_ ( .D(n10520), .CLK(clk), .Q(arr[2218]) );
  DFFPOSX1 arr_reg_54__3_ ( .D(n10519), .CLK(clk), .Q(arr[2217]) );
  DFFPOSX1 arr_reg_54__2_ ( .D(n10518), .CLK(clk), .Q(arr[2216]) );
  DFFPOSX1 arr_reg_54__1_ ( .D(n10517), .CLK(clk), .Q(arr[2215]) );
  DFFPOSX1 arr_reg_54__0_ ( .D(n10516), .CLK(clk), .Q(arr[2214]) );
  DFFPOSX1 arr_reg_53__40_ ( .D(n10515), .CLK(clk), .Q(arr[2213]) );
  DFFPOSX1 arr_reg_53__39_ ( .D(n10514), .CLK(clk), .Q(arr[2212]) );
  DFFPOSX1 arr_reg_53__38_ ( .D(n10513), .CLK(clk), .Q(arr[2211]) );
  DFFPOSX1 arr_reg_53__37_ ( .D(n10512), .CLK(clk), .Q(arr[2210]) );
  DFFPOSX1 arr_reg_53__36_ ( .D(n10511), .CLK(clk), .Q(arr[2209]) );
  DFFPOSX1 arr_reg_53__35_ ( .D(n10510), .CLK(clk), .Q(arr[2208]) );
  DFFPOSX1 arr_reg_53__34_ ( .D(n10509), .CLK(clk), .Q(arr[2207]) );
  DFFPOSX1 arr_reg_53__33_ ( .D(n10508), .CLK(clk), .Q(arr[2206]) );
  DFFPOSX1 arr_reg_53__32_ ( .D(n10507), .CLK(clk), .Q(arr[2205]) );
  DFFPOSX1 arr_reg_53__31_ ( .D(n10506), .CLK(clk), .Q(arr[2204]) );
  DFFPOSX1 arr_reg_53__30_ ( .D(n10505), .CLK(clk), .Q(arr[2203]) );
  DFFPOSX1 arr_reg_53__29_ ( .D(n10504), .CLK(clk), .Q(arr[2202]) );
  DFFPOSX1 arr_reg_53__28_ ( .D(n10503), .CLK(clk), .Q(arr[2201]) );
  DFFPOSX1 arr_reg_53__27_ ( .D(n10502), .CLK(clk), .Q(arr[2200]) );
  DFFPOSX1 arr_reg_53__26_ ( .D(n10501), .CLK(clk), .Q(arr[2199]) );
  DFFPOSX1 arr_reg_53__25_ ( .D(n10500), .CLK(clk), .Q(arr[2198]) );
  DFFPOSX1 arr_reg_53__24_ ( .D(n10499), .CLK(clk), .Q(arr[2197]) );
  DFFPOSX1 arr_reg_53__23_ ( .D(n10498), .CLK(clk), .Q(arr[2196]) );
  DFFPOSX1 arr_reg_53__22_ ( .D(n10497), .CLK(clk), .Q(arr[2195]) );
  DFFPOSX1 arr_reg_53__21_ ( .D(n10496), .CLK(clk), .Q(arr[2194]) );
  DFFPOSX1 arr_reg_53__20_ ( .D(n10495), .CLK(clk), .Q(arr[2193]) );
  DFFPOSX1 arr_reg_53__19_ ( .D(n10494), .CLK(clk), .Q(arr[2192]) );
  DFFPOSX1 arr_reg_53__18_ ( .D(n10493), .CLK(clk), .Q(arr[2191]) );
  DFFPOSX1 arr_reg_53__17_ ( .D(n10492), .CLK(clk), .Q(arr[2190]) );
  DFFPOSX1 arr_reg_53__16_ ( .D(n10491), .CLK(clk), .Q(arr[2189]) );
  DFFPOSX1 arr_reg_53__15_ ( .D(n10490), .CLK(clk), .Q(arr[2188]) );
  DFFPOSX1 arr_reg_53__14_ ( .D(n10489), .CLK(clk), .Q(arr[2187]) );
  DFFPOSX1 arr_reg_53__13_ ( .D(n10488), .CLK(clk), .Q(arr[2186]) );
  DFFPOSX1 arr_reg_53__12_ ( .D(n10487), .CLK(clk), .Q(arr[2185]) );
  DFFPOSX1 arr_reg_53__11_ ( .D(n10486), .CLK(clk), .Q(arr[2184]) );
  DFFPOSX1 arr_reg_53__10_ ( .D(n10485), .CLK(clk), .Q(arr[2183]) );
  DFFPOSX1 arr_reg_53__9_ ( .D(n10484), .CLK(clk), .Q(arr[2182]) );
  DFFPOSX1 arr_reg_53__8_ ( .D(n10483), .CLK(clk), .Q(arr[2181]) );
  DFFPOSX1 arr_reg_53__7_ ( .D(n10482), .CLK(clk), .Q(arr[2180]) );
  DFFPOSX1 arr_reg_53__6_ ( .D(n10481), .CLK(clk), .Q(arr[2179]) );
  DFFPOSX1 arr_reg_53__5_ ( .D(n10480), .CLK(clk), .Q(arr[2178]) );
  DFFPOSX1 arr_reg_53__4_ ( .D(n10479), .CLK(clk), .Q(arr[2177]) );
  DFFPOSX1 arr_reg_53__3_ ( .D(n10478), .CLK(clk), .Q(arr[2176]) );
  DFFPOSX1 arr_reg_53__2_ ( .D(n10477), .CLK(clk), .Q(arr[2175]) );
  DFFPOSX1 arr_reg_53__1_ ( .D(n10476), .CLK(clk), .Q(arr[2174]) );
  DFFPOSX1 arr_reg_53__0_ ( .D(n10475), .CLK(clk), .Q(arr[2173]) );
  DFFPOSX1 arr_reg_52__40_ ( .D(n10474), .CLK(clk), .Q(arr[2172]) );
  DFFPOSX1 arr_reg_52__39_ ( .D(n10473), .CLK(clk), .Q(arr[2171]) );
  DFFPOSX1 arr_reg_52__38_ ( .D(n10472), .CLK(clk), .Q(arr[2170]) );
  DFFPOSX1 arr_reg_52__37_ ( .D(n10471), .CLK(clk), .Q(arr[2169]) );
  DFFPOSX1 arr_reg_52__36_ ( .D(n10470), .CLK(clk), .Q(arr[2168]) );
  DFFPOSX1 arr_reg_52__35_ ( .D(n10469), .CLK(clk), .Q(arr[2167]) );
  DFFPOSX1 arr_reg_52__34_ ( .D(n10468), .CLK(clk), .Q(arr[2166]) );
  DFFPOSX1 arr_reg_52__33_ ( .D(n10467), .CLK(clk), .Q(arr[2165]) );
  DFFPOSX1 arr_reg_52__32_ ( .D(n10466), .CLK(clk), .Q(arr[2164]) );
  DFFPOSX1 arr_reg_52__31_ ( .D(n10465), .CLK(clk), .Q(arr[2163]) );
  DFFPOSX1 arr_reg_52__30_ ( .D(n10464), .CLK(clk), .Q(arr[2162]) );
  DFFPOSX1 arr_reg_52__29_ ( .D(n10463), .CLK(clk), .Q(arr[2161]) );
  DFFPOSX1 arr_reg_52__28_ ( .D(n10462), .CLK(clk), .Q(arr[2160]) );
  DFFPOSX1 arr_reg_52__27_ ( .D(n10461), .CLK(clk), .Q(arr[2159]) );
  DFFPOSX1 arr_reg_52__26_ ( .D(n10460), .CLK(clk), .Q(arr[2158]) );
  DFFPOSX1 arr_reg_52__25_ ( .D(n10459), .CLK(clk), .Q(arr[2157]) );
  DFFPOSX1 arr_reg_52__24_ ( .D(n10458), .CLK(clk), .Q(arr[2156]) );
  DFFPOSX1 arr_reg_52__23_ ( .D(n10457), .CLK(clk), .Q(arr[2155]) );
  DFFPOSX1 arr_reg_52__22_ ( .D(n10456), .CLK(clk), .Q(arr[2154]) );
  DFFPOSX1 arr_reg_52__21_ ( .D(n10455), .CLK(clk), .Q(arr[2153]) );
  DFFPOSX1 arr_reg_52__20_ ( .D(n10454), .CLK(clk), .Q(arr[2152]) );
  DFFPOSX1 arr_reg_52__19_ ( .D(n10453), .CLK(clk), .Q(arr[2151]) );
  DFFPOSX1 arr_reg_52__18_ ( .D(n10452), .CLK(clk), .Q(arr[2150]) );
  DFFPOSX1 arr_reg_52__17_ ( .D(n10451), .CLK(clk), .Q(arr[2149]) );
  DFFPOSX1 arr_reg_52__16_ ( .D(n10450), .CLK(clk), .Q(arr[2148]) );
  DFFPOSX1 arr_reg_52__15_ ( .D(n10449), .CLK(clk), .Q(arr[2147]) );
  DFFPOSX1 arr_reg_52__14_ ( .D(n10448), .CLK(clk), .Q(arr[2146]) );
  DFFPOSX1 arr_reg_52__13_ ( .D(n10447), .CLK(clk), .Q(arr[2145]) );
  DFFPOSX1 arr_reg_52__12_ ( .D(n10446), .CLK(clk), .Q(arr[2144]) );
  DFFPOSX1 arr_reg_52__11_ ( .D(n10445), .CLK(clk), .Q(arr[2143]) );
  DFFPOSX1 arr_reg_52__10_ ( .D(n10444), .CLK(clk), .Q(arr[2142]) );
  DFFPOSX1 arr_reg_52__9_ ( .D(n10443), .CLK(clk), .Q(arr[2141]) );
  DFFPOSX1 arr_reg_52__8_ ( .D(n10442), .CLK(clk), .Q(arr[2140]) );
  DFFPOSX1 arr_reg_52__7_ ( .D(n10441), .CLK(clk), .Q(arr[2139]) );
  DFFPOSX1 arr_reg_52__6_ ( .D(n10440), .CLK(clk), .Q(arr[2138]) );
  DFFPOSX1 arr_reg_52__5_ ( .D(n10439), .CLK(clk), .Q(arr[2137]) );
  DFFPOSX1 arr_reg_52__4_ ( .D(n10438), .CLK(clk), .Q(arr[2136]) );
  DFFPOSX1 arr_reg_52__3_ ( .D(n10437), .CLK(clk), .Q(arr[2135]) );
  DFFPOSX1 arr_reg_52__2_ ( .D(n10436), .CLK(clk), .Q(arr[2134]) );
  DFFPOSX1 arr_reg_52__1_ ( .D(n10435), .CLK(clk), .Q(arr[2133]) );
  DFFPOSX1 arr_reg_52__0_ ( .D(n10434), .CLK(clk), .Q(arr[2132]) );
  DFFPOSX1 arr_reg_51__40_ ( .D(n10433), .CLK(clk), .Q(arr[2131]) );
  DFFPOSX1 arr_reg_51__39_ ( .D(n10432), .CLK(clk), .Q(arr[2130]) );
  DFFPOSX1 arr_reg_51__38_ ( .D(n10431), .CLK(clk), .Q(arr[2129]) );
  DFFPOSX1 arr_reg_51__37_ ( .D(n10430), .CLK(clk), .Q(arr[2128]) );
  DFFPOSX1 arr_reg_51__36_ ( .D(n10429), .CLK(clk), .Q(arr[2127]) );
  DFFPOSX1 arr_reg_51__35_ ( .D(n10428), .CLK(clk), .Q(arr[2126]) );
  DFFPOSX1 arr_reg_51__34_ ( .D(n10427), .CLK(clk), .Q(arr[2125]) );
  DFFPOSX1 arr_reg_51__33_ ( .D(n10426), .CLK(clk), .Q(arr[2124]) );
  DFFPOSX1 arr_reg_51__32_ ( .D(n10425), .CLK(clk), .Q(arr[2123]) );
  DFFPOSX1 arr_reg_51__31_ ( .D(n10424), .CLK(clk), .Q(arr[2122]) );
  DFFPOSX1 arr_reg_51__30_ ( .D(n10423), .CLK(clk), .Q(arr[2121]) );
  DFFPOSX1 arr_reg_51__29_ ( .D(n10422), .CLK(clk), .Q(arr[2120]) );
  DFFPOSX1 arr_reg_51__28_ ( .D(n10421), .CLK(clk), .Q(arr[2119]) );
  DFFPOSX1 arr_reg_51__27_ ( .D(n10420), .CLK(clk), .Q(arr[2118]) );
  DFFPOSX1 arr_reg_51__26_ ( .D(n10419), .CLK(clk), .Q(arr[2117]) );
  DFFPOSX1 arr_reg_51__25_ ( .D(n10418), .CLK(clk), .Q(arr[2116]) );
  DFFPOSX1 arr_reg_51__24_ ( .D(n10417), .CLK(clk), .Q(arr[2115]) );
  DFFPOSX1 arr_reg_51__23_ ( .D(n10416), .CLK(clk), .Q(arr[2114]) );
  DFFPOSX1 arr_reg_51__22_ ( .D(n10415), .CLK(clk), .Q(arr[2113]) );
  DFFPOSX1 arr_reg_51__21_ ( .D(n10414), .CLK(clk), .Q(arr[2112]) );
  DFFPOSX1 arr_reg_51__20_ ( .D(n10413), .CLK(clk), .Q(arr[2111]) );
  DFFPOSX1 arr_reg_51__19_ ( .D(n10412), .CLK(clk), .Q(arr[2110]) );
  DFFPOSX1 arr_reg_51__18_ ( .D(n10411), .CLK(clk), .Q(arr[2109]) );
  DFFPOSX1 arr_reg_51__17_ ( .D(n10410), .CLK(clk), .Q(arr[2108]) );
  DFFPOSX1 arr_reg_51__16_ ( .D(n10409), .CLK(clk), .Q(arr[2107]) );
  DFFPOSX1 arr_reg_51__15_ ( .D(n10408), .CLK(clk), .Q(arr[2106]) );
  DFFPOSX1 arr_reg_51__14_ ( .D(n10407), .CLK(clk), .Q(arr[2105]) );
  DFFPOSX1 arr_reg_51__13_ ( .D(n10406), .CLK(clk), .Q(arr[2104]) );
  DFFPOSX1 arr_reg_51__12_ ( .D(n10405), .CLK(clk), .Q(arr[2103]) );
  DFFPOSX1 arr_reg_51__11_ ( .D(n10404), .CLK(clk), .Q(arr[2102]) );
  DFFPOSX1 arr_reg_51__10_ ( .D(n10403), .CLK(clk), .Q(arr[2101]) );
  DFFPOSX1 arr_reg_51__9_ ( .D(n10402), .CLK(clk), .Q(arr[2100]) );
  DFFPOSX1 arr_reg_51__8_ ( .D(n10401), .CLK(clk), .Q(arr[2099]) );
  DFFPOSX1 arr_reg_51__7_ ( .D(n10400), .CLK(clk), .Q(arr[2098]) );
  DFFPOSX1 arr_reg_51__6_ ( .D(n10399), .CLK(clk), .Q(arr[2097]) );
  DFFPOSX1 arr_reg_51__5_ ( .D(n10398), .CLK(clk), .Q(arr[2096]) );
  DFFPOSX1 arr_reg_51__4_ ( .D(n10397), .CLK(clk), .Q(arr[2095]) );
  DFFPOSX1 arr_reg_51__3_ ( .D(n10396), .CLK(clk), .Q(arr[2094]) );
  DFFPOSX1 arr_reg_51__2_ ( .D(n10395), .CLK(clk), .Q(arr[2093]) );
  DFFPOSX1 arr_reg_51__1_ ( .D(n10394), .CLK(clk), .Q(arr[2092]) );
  DFFPOSX1 arr_reg_51__0_ ( .D(n10393), .CLK(clk), .Q(arr[2091]) );
  DFFPOSX1 arr_reg_50__40_ ( .D(n10392), .CLK(clk), .Q(arr[2090]) );
  DFFPOSX1 arr_reg_50__39_ ( .D(n10391), .CLK(clk), .Q(arr[2089]) );
  DFFPOSX1 arr_reg_50__38_ ( .D(n10390), .CLK(clk), .Q(arr[2088]) );
  DFFPOSX1 arr_reg_50__37_ ( .D(n10389), .CLK(clk), .Q(arr[2087]) );
  DFFPOSX1 arr_reg_50__36_ ( .D(n10388), .CLK(clk), .Q(arr[2086]) );
  DFFPOSX1 arr_reg_50__35_ ( .D(n10387), .CLK(clk), .Q(arr[2085]) );
  DFFPOSX1 arr_reg_50__34_ ( .D(n10386), .CLK(clk), .Q(arr[2084]) );
  DFFPOSX1 arr_reg_50__33_ ( .D(n10385), .CLK(clk), .Q(arr[2083]) );
  DFFPOSX1 arr_reg_50__32_ ( .D(n10384), .CLK(clk), .Q(arr[2082]) );
  DFFPOSX1 arr_reg_50__31_ ( .D(n10383), .CLK(clk), .Q(arr[2081]) );
  DFFPOSX1 arr_reg_50__30_ ( .D(n10382), .CLK(clk), .Q(arr[2080]) );
  DFFPOSX1 arr_reg_50__29_ ( .D(n10381), .CLK(clk), .Q(arr[2079]) );
  DFFPOSX1 arr_reg_50__28_ ( .D(n10380), .CLK(clk), .Q(arr[2078]) );
  DFFPOSX1 arr_reg_50__27_ ( .D(n10379), .CLK(clk), .Q(arr[2077]) );
  DFFPOSX1 arr_reg_50__26_ ( .D(n10378), .CLK(clk), .Q(arr[2076]) );
  DFFPOSX1 arr_reg_50__25_ ( .D(n10377), .CLK(clk), .Q(arr[2075]) );
  DFFPOSX1 arr_reg_50__24_ ( .D(n10376), .CLK(clk), .Q(arr[2074]) );
  DFFPOSX1 arr_reg_50__23_ ( .D(n10375), .CLK(clk), .Q(arr[2073]) );
  DFFPOSX1 arr_reg_50__22_ ( .D(n10374), .CLK(clk), .Q(arr[2072]) );
  DFFPOSX1 arr_reg_50__21_ ( .D(n10373), .CLK(clk), .Q(arr[2071]) );
  DFFPOSX1 arr_reg_50__20_ ( .D(n10372), .CLK(clk), .Q(arr[2070]) );
  DFFPOSX1 arr_reg_50__19_ ( .D(n10371), .CLK(clk), .Q(arr[2069]) );
  DFFPOSX1 arr_reg_50__18_ ( .D(n10370), .CLK(clk), .Q(arr[2068]) );
  DFFPOSX1 arr_reg_50__17_ ( .D(n10369), .CLK(clk), .Q(arr[2067]) );
  DFFPOSX1 arr_reg_50__16_ ( .D(n10368), .CLK(clk), .Q(arr[2066]) );
  DFFPOSX1 arr_reg_50__15_ ( .D(n10367), .CLK(clk), .Q(arr[2065]) );
  DFFPOSX1 arr_reg_50__14_ ( .D(n10366), .CLK(clk), .Q(arr[2064]) );
  DFFPOSX1 arr_reg_50__13_ ( .D(n10365), .CLK(clk), .Q(arr[2063]) );
  DFFPOSX1 arr_reg_50__12_ ( .D(n10364), .CLK(clk), .Q(arr[2062]) );
  DFFPOSX1 arr_reg_50__11_ ( .D(n10363), .CLK(clk), .Q(arr[2061]) );
  DFFPOSX1 arr_reg_50__10_ ( .D(n10362), .CLK(clk), .Q(arr[2060]) );
  DFFPOSX1 arr_reg_50__9_ ( .D(n10361), .CLK(clk), .Q(arr[2059]) );
  DFFPOSX1 arr_reg_50__8_ ( .D(n10360), .CLK(clk), .Q(arr[2058]) );
  DFFPOSX1 arr_reg_50__7_ ( .D(n10359), .CLK(clk), .Q(arr[2057]) );
  DFFPOSX1 arr_reg_50__6_ ( .D(n10358), .CLK(clk), .Q(arr[2056]) );
  DFFPOSX1 arr_reg_50__5_ ( .D(n10357), .CLK(clk), .Q(arr[2055]) );
  DFFPOSX1 arr_reg_50__4_ ( .D(n10356), .CLK(clk), .Q(arr[2054]) );
  DFFPOSX1 arr_reg_50__3_ ( .D(n10355), .CLK(clk), .Q(arr[2053]) );
  DFFPOSX1 arr_reg_50__2_ ( .D(n10354), .CLK(clk), .Q(arr[2052]) );
  DFFPOSX1 arr_reg_50__1_ ( .D(n10353), .CLK(clk), .Q(arr[2051]) );
  DFFPOSX1 arr_reg_50__0_ ( .D(n10352), .CLK(clk), .Q(arr[2050]) );
  DFFPOSX1 arr_reg_49__40_ ( .D(n10351), .CLK(clk), .Q(arr[2049]) );
  DFFPOSX1 arr_reg_49__39_ ( .D(n10350), .CLK(clk), .Q(arr[2048]) );
  DFFPOSX1 arr_reg_49__38_ ( .D(n10349), .CLK(clk), .Q(arr[2047]) );
  DFFPOSX1 arr_reg_49__37_ ( .D(n10348), .CLK(clk), .Q(arr[2046]) );
  DFFPOSX1 arr_reg_49__36_ ( .D(n10347), .CLK(clk), .Q(arr[2045]) );
  DFFPOSX1 arr_reg_49__35_ ( .D(n10346), .CLK(clk), .Q(arr[2044]) );
  DFFPOSX1 arr_reg_49__34_ ( .D(n10345), .CLK(clk), .Q(arr[2043]) );
  DFFPOSX1 arr_reg_49__33_ ( .D(n10344), .CLK(clk), .Q(arr[2042]) );
  DFFPOSX1 arr_reg_49__32_ ( .D(n10343), .CLK(clk), .Q(arr[2041]) );
  DFFPOSX1 arr_reg_49__31_ ( .D(n10342), .CLK(clk), .Q(arr[2040]) );
  DFFPOSX1 arr_reg_49__30_ ( .D(n10341), .CLK(clk), .Q(arr[2039]) );
  DFFPOSX1 arr_reg_49__29_ ( .D(n10340), .CLK(clk), .Q(arr[2038]) );
  DFFPOSX1 arr_reg_49__28_ ( .D(n10339), .CLK(clk), .Q(arr[2037]) );
  DFFPOSX1 arr_reg_49__27_ ( .D(n10338), .CLK(clk), .Q(arr[2036]) );
  DFFPOSX1 arr_reg_49__26_ ( .D(n10337), .CLK(clk), .Q(arr[2035]) );
  DFFPOSX1 arr_reg_49__25_ ( .D(n10336), .CLK(clk), .Q(arr[2034]) );
  DFFPOSX1 arr_reg_49__24_ ( .D(n10335), .CLK(clk), .Q(arr[2033]) );
  DFFPOSX1 arr_reg_49__23_ ( .D(n10334), .CLK(clk), .Q(arr[2032]) );
  DFFPOSX1 arr_reg_49__22_ ( .D(n10333), .CLK(clk), .Q(arr[2031]) );
  DFFPOSX1 arr_reg_49__21_ ( .D(n10332), .CLK(clk), .Q(arr[2030]) );
  DFFPOSX1 arr_reg_49__20_ ( .D(n10331), .CLK(clk), .Q(arr[2029]) );
  DFFPOSX1 arr_reg_49__19_ ( .D(n10330), .CLK(clk), .Q(arr[2028]) );
  DFFPOSX1 arr_reg_49__18_ ( .D(n10329), .CLK(clk), .Q(arr[2027]) );
  DFFPOSX1 arr_reg_49__17_ ( .D(n10328), .CLK(clk), .Q(arr[2026]) );
  DFFPOSX1 arr_reg_49__16_ ( .D(n10327), .CLK(clk), .Q(arr[2025]) );
  DFFPOSX1 arr_reg_49__15_ ( .D(n10326), .CLK(clk), .Q(arr[2024]) );
  DFFPOSX1 arr_reg_49__14_ ( .D(n10325), .CLK(clk), .Q(arr[2023]) );
  DFFPOSX1 arr_reg_49__13_ ( .D(n10324), .CLK(clk), .Q(arr[2022]) );
  DFFPOSX1 arr_reg_49__12_ ( .D(n10323), .CLK(clk), .Q(arr[2021]) );
  DFFPOSX1 arr_reg_49__11_ ( .D(n10322), .CLK(clk), .Q(arr[2020]) );
  DFFPOSX1 arr_reg_49__10_ ( .D(n10321), .CLK(clk), .Q(arr[2019]) );
  DFFPOSX1 arr_reg_49__9_ ( .D(n10320), .CLK(clk), .Q(arr[2018]) );
  DFFPOSX1 arr_reg_49__8_ ( .D(n10319), .CLK(clk), .Q(arr[2017]) );
  DFFPOSX1 arr_reg_49__7_ ( .D(n10318), .CLK(clk), .Q(arr[2016]) );
  DFFPOSX1 arr_reg_49__6_ ( .D(n10317), .CLK(clk), .Q(arr[2015]) );
  DFFPOSX1 arr_reg_49__5_ ( .D(n10316), .CLK(clk), .Q(arr[2014]) );
  DFFPOSX1 arr_reg_49__4_ ( .D(n10315), .CLK(clk), .Q(arr[2013]) );
  DFFPOSX1 arr_reg_49__3_ ( .D(n10314), .CLK(clk), .Q(arr[2012]) );
  DFFPOSX1 arr_reg_49__2_ ( .D(n10313), .CLK(clk), .Q(arr[2011]) );
  DFFPOSX1 arr_reg_49__1_ ( .D(n10312), .CLK(clk), .Q(arr[2010]) );
  DFFPOSX1 arr_reg_49__0_ ( .D(n10311), .CLK(clk), .Q(arr[2009]) );
  DFFPOSX1 arr_reg_48__40_ ( .D(n10310), .CLK(clk), .Q(arr[2008]) );
  DFFPOSX1 arr_reg_48__39_ ( .D(n10309), .CLK(clk), .Q(arr[2007]) );
  DFFPOSX1 arr_reg_48__38_ ( .D(n10308), .CLK(clk), .Q(arr[2006]) );
  DFFPOSX1 arr_reg_48__37_ ( .D(n10307), .CLK(clk), .Q(arr[2005]) );
  DFFPOSX1 arr_reg_48__36_ ( .D(n10306), .CLK(clk), .Q(arr[2004]) );
  DFFPOSX1 arr_reg_48__35_ ( .D(n10305), .CLK(clk), .Q(arr[2003]) );
  DFFPOSX1 arr_reg_48__34_ ( .D(n10304), .CLK(clk), .Q(arr[2002]) );
  DFFPOSX1 arr_reg_48__33_ ( .D(n10303), .CLK(clk), .Q(arr[2001]) );
  DFFPOSX1 arr_reg_48__32_ ( .D(n10302), .CLK(clk), .Q(arr[2000]) );
  DFFPOSX1 arr_reg_48__31_ ( .D(n10301), .CLK(clk), .Q(arr[1999]) );
  DFFPOSX1 arr_reg_48__30_ ( .D(n10300), .CLK(clk), .Q(arr[1998]) );
  DFFPOSX1 arr_reg_48__29_ ( .D(n10299), .CLK(clk), .Q(arr[1997]) );
  DFFPOSX1 arr_reg_48__28_ ( .D(n10298), .CLK(clk), .Q(arr[1996]) );
  DFFPOSX1 arr_reg_48__27_ ( .D(n10297), .CLK(clk), .Q(arr[1995]) );
  DFFPOSX1 arr_reg_48__26_ ( .D(n10296), .CLK(clk), .Q(arr[1994]) );
  DFFPOSX1 arr_reg_48__25_ ( .D(n10295), .CLK(clk), .Q(arr[1993]) );
  DFFPOSX1 arr_reg_48__24_ ( .D(n10294), .CLK(clk), .Q(arr[1992]) );
  DFFPOSX1 arr_reg_48__23_ ( .D(n10293), .CLK(clk), .Q(arr[1991]) );
  DFFPOSX1 arr_reg_48__22_ ( .D(n10292), .CLK(clk), .Q(arr[1990]) );
  DFFPOSX1 arr_reg_48__21_ ( .D(n10291), .CLK(clk), .Q(arr[1989]) );
  DFFPOSX1 arr_reg_48__20_ ( .D(n10290), .CLK(clk), .Q(arr[1988]) );
  DFFPOSX1 arr_reg_48__19_ ( .D(n10289), .CLK(clk), .Q(arr[1987]) );
  DFFPOSX1 arr_reg_48__18_ ( .D(n10288), .CLK(clk), .Q(arr[1986]) );
  DFFPOSX1 arr_reg_48__17_ ( .D(n10287), .CLK(clk), .Q(arr[1985]) );
  DFFPOSX1 arr_reg_48__16_ ( .D(n10286), .CLK(clk), .Q(arr[1984]) );
  DFFPOSX1 arr_reg_48__15_ ( .D(n10285), .CLK(clk), .Q(arr[1983]) );
  DFFPOSX1 arr_reg_48__14_ ( .D(n10284), .CLK(clk), .Q(arr[1982]) );
  DFFPOSX1 arr_reg_48__13_ ( .D(n10283), .CLK(clk), .Q(arr[1981]) );
  DFFPOSX1 arr_reg_48__12_ ( .D(n10282), .CLK(clk), .Q(arr[1980]) );
  DFFPOSX1 arr_reg_48__11_ ( .D(n10281), .CLK(clk), .Q(arr[1979]) );
  DFFPOSX1 arr_reg_48__10_ ( .D(n10280), .CLK(clk), .Q(arr[1978]) );
  DFFPOSX1 arr_reg_48__9_ ( .D(n10279), .CLK(clk), .Q(arr[1977]) );
  DFFPOSX1 arr_reg_48__8_ ( .D(n10278), .CLK(clk), .Q(arr[1976]) );
  DFFPOSX1 arr_reg_48__7_ ( .D(n10277), .CLK(clk), .Q(arr[1975]) );
  DFFPOSX1 arr_reg_48__6_ ( .D(n10276), .CLK(clk), .Q(arr[1974]) );
  DFFPOSX1 arr_reg_48__5_ ( .D(n10275), .CLK(clk), .Q(arr[1973]) );
  DFFPOSX1 arr_reg_48__4_ ( .D(n10274), .CLK(clk), .Q(arr[1972]) );
  DFFPOSX1 arr_reg_48__3_ ( .D(n10273), .CLK(clk), .Q(arr[1971]) );
  DFFPOSX1 arr_reg_48__2_ ( .D(n10272), .CLK(clk), .Q(arr[1970]) );
  DFFPOSX1 arr_reg_48__1_ ( .D(n10271), .CLK(clk), .Q(arr[1969]) );
  DFFPOSX1 arr_reg_48__0_ ( .D(n10270), .CLK(clk), .Q(arr[1968]) );
  DFFPOSX1 arr_reg_47__40_ ( .D(n10269), .CLK(clk), .Q(arr[1967]) );
  DFFPOSX1 arr_reg_47__39_ ( .D(n10268), .CLK(clk), .Q(arr[1966]) );
  DFFPOSX1 arr_reg_47__38_ ( .D(n10267), .CLK(clk), .Q(arr[1965]) );
  DFFPOSX1 arr_reg_47__37_ ( .D(n10266), .CLK(clk), .Q(arr[1964]) );
  DFFPOSX1 arr_reg_47__36_ ( .D(n10265), .CLK(clk), .Q(arr[1963]) );
  DFFPOSX1 arr_reg_47__35_ ( .D(n10264), .CLK(clk), .Q(arr[1962]) );
  DFFPOSX1 arr_reg_47__34_ ( .D(n10263), .CLK(clk), .Q(arr[1961]) );
  DFFPOSX1 arr_reg_47__33_ ( .D(n10262), .CLK(clk), .Q(arr[1960]) );
  DFFPOSX1 arr_reg_47__32_ ( .D(n10261), .CLK(clk), .Q(arr[1959]) );
  DFFPOSX1 arr_reg_47__31_ ( .D(n10260), .CLK(clk), .Q(arr[1958]) );
  DFFPOSX1 arr_reg_47__30_ ( .D(n10259), .CLK(clk), .Q(arr[1957]) );
  DFFPOSX1 arr_reg_47__29_ ( .D(n10258), .CLK(clk), .Q(arr[1956]) );
  DFFPOSX1 arr_reg_47__28_ ( .D(n10257), .CLK(clk), .Q(arr[1955]) );
  DFFPOSX1 arr_reg_47__27_ ( .D(n10256), .CLK(clk), .Q(arr[1954]) );
  DFFPOSX1 arr_reg_47__26_ ( .D(n10255), .CLK(clk), .Q(arr[1953]) );
  DFFPOSX1 arr_reg_47__25_ ( .D(n10254), .CLK(clk), .Q(arr[1952]) );
  DFFPOSX1 arr_reg_47__24_ ( .D(n10253), .CLK(clk), .Q(arr[1951]) );
  DFFPOSX1 arr_reg_47__23_ ( .D(n10252), .CLK(clk), .Q(arr[1950]) );
  DFFPOSX1 arr_reg_47__22_ ( .D(n10251), .CLK(clk), .Q(arr[1949]) );
  DFFPOSX1 arr_reg_47__21_ ( .D(n10250), .CLK(clk), .Q(arr[1948]) );
  DFFPOSX1 arr_reg_47__20_ ( .D(n10249), .CLK(clk), .Q(arr[1947]) );
  DFFPOSX1 arr_reg_47__19_ ( .D(n10248), .CLK(clk), .Q(arr[1946]) );
  DFFPOSX1 arr_reg_47__18_ ( .D(n10247), .CLK(clk), .Q(arr[1945]) );
  DFFPOSX1 arr_reg_47__17_ ( .D(n10246), .CLK(clk), .Q(arr[1944]) );
  DFFPOSX1 arr_reg_47__16_ ( .D(n10245), .CLK(clk), .Q(arr[1943]) );
  DFFPOSX1 arr_reg_47__15_ ( .D(n10244), .CLK(clk), .Q(arr[1942]) );
  DFFPOSX1 arr_reg_47__14_ ( .D(n10243), .CLK(clk), .Q(arr[1941]) );
  DFFPOSX1 arr_reg_47__13_ ( .D(n10242), .CLK(clk), .Q(arr[1940]) );
  DFFPOSX1 arr_reg_47__12_ ( .D(n10241), .CLK(clk), .Q(arr[1939]) );
  DFFPOSX1 arr_reg_47__11_ ( .D(n10240), .CLK(clk), .Q(arr[1938]) );
  DFFPOSX1 arr_reg_47__10_ ( .D(n10239), .CLK(clk), .Q(arr[1937]) );
  DFFPOSX1 arr_reg_47__9_ ( .D(n10238), .CLK(clk), .Q(arr[1936]) );
  DFFPOSX1 arr_reg_47__8_ ( .D(n10237), .CLK(clk), .Q(arr[1935]) );
  DFFPOSX1 arr_reg_47__7_ ( .D(n10236), .CLK(clk), .Q(arr[1934]) );
  DFFPOSX1 arr_reg_47__6_ ( .D(n10235), .CLK(clk), .Q(arr[1933]) );
  DFFPOSX1 arr_reg_47__5_ ( .D(n10234), .CLK(clk), .Q(arr[1932]) );
  DFFPOSX1 arr_reg_47__4_ ( .D(n10233), .CLK(clk), .Q(arr[1931]) );
  DFFPOSX1 arr_reg_47__3_ ( .D(n10232), .CLK(clk), .Q(arr[1930]) );
  DFFPOSX1 arr_reg_47__2_ ( .D(n10231), .CLK(clk), .Q(arr[1929]) );
  DFFPOSX1 arr_reg_47__1_ ( .D(n10230), .CLK(clk), .Q(arr[1928]) );
  DFFPOSX1 arr_reg_47__0_ ( .D(n10229), .CLK(clk), .Q(arr[1927]) );
  DFFPOSX1 arr_reg_46__40_ ( .D(n10228), .CLK(clk), .Q(arr[1926]) );
  DFFPOSX1 arr_reg_46__39_ ( .D(n10227), .CLK(clk), .Q(arr[1925]) );
  DFFPOSX1 arr_reg_46__38_ ( .D(n10226), .CLK(clk), .Q(arr[1924]) );
  DFFPOSX1 arr_reg_46__37_ ( .D(n10225), .CLK(clk), .Q(arr[1923]) );
  DFFPOSX1 arr_reg_46__36_ ( .D(n10224), .CLK(clk), .Q(arr[1922]) );
  DFFPOSX1 arr_reg_46__35_ ( .D(n10223), .CLK(clk), .Q(arr[1921]) );
  DFFPOSX1 arr_reg_46__34_ ( .D(n10222), .CLK(clk), .Q(arr[1920]) );
  DFFPOSX1 arr_reg_46__33_ ( .D(n10221), .CLK(clk), .Q(arr[1919]) );
  DFFPOSX1 arr_reg_46__32_ ( .D(n10220), .CLK(clk), .Q(arr[1918]) );
  DFFPOSX1 arr_reg_46__31_ ( .D(n10219), .CLK(clk), .Q(arr[1917]) );
  DFFPOSX1 arr_reg_46__30_ ( .D(n10218), .CLK(clk), .Q(arr[1916]) );
  DFFPOSX1 arr_reg_46__29_ ( .D(n10217), .CLK(clk), .Q(arr[1915]) );
  DFFPOSX1 arr_reg_46__28_ ( .D(n10216), .CLK(clk), .Q(arr[1914]) );
  DFFPOSX1 arr_reg_46__27_ ( .D(n10215), .CLK(clk), .Q(arr[1913]) );
  DFFPOSX1 arr_reg_46__26_ ( .D(n10214), .CLK(clk), .Q(arr[1912]) );
  DFFPOSX1 arr_reg_46__25_ ( .D(n10213), .CLK(clk), .Q(arr[1911]) );
  DFFPOSX1 arr_reg_46__24_ ( .D(n10212), .CLK(clk), .Q(arr[1910]) );
  DFFPOSX1 arr_reg_46__23_ ( .D(n10211), .CLK(clk), .Q(arr[1909]) );
  DFFPOSX1 arr_reg_46__22_ ( .D(n10210), .CLK(clk), .Q(arr[1908]) );
  DFFPOSX1 arr_reg_46__21_ ( .D(n10209), .CLK(clk), .Q(arr[1907]) );
  DFFPOSX1 arr_reg_46__20_ ( .D(n10208), .CLK(clk), .Q(arr[1906]) );
  DFFPOSX1 arr_reg_46__19_ ( .D(n10207), .CLK(clk), .Q(arr[1905]) );
  DFFPOSX1 arr_reg_46__18_ ( .D(n10206), .CLK(clk), .Q(arr[1904]) );
  DFFPOSX1 arr_reg_46__17_ ( .D(n10205), .CLK(clk), .Q(arr[1903]) );
  DFFPOSX1 arr_reg_46__16_ ( .D(n10204), .CLK(clk), .Q(arr[1902]) );
  DFFPOSX1 arr_reg_46__15_ ( .D(n10203), .CLK(clk), .Q(arr[1901]) );
  DFFPOSX1 arr_reg_46__14_ ( .D(n10202), .CLK(clk), .Q(arr[1900]) );
  DFFPOSX1 arr_reg_46__13_ ( .D(n10201), .CLK(clk), .Q(arr[1899]) );
  DFFPOSX1 arr_reg_46__12_ ( .D(n10200), .CLK(clk), .Q(arr[1898]) );
  DFFPOSX1 arr_reg_46__11_ ( .D(n10199), .CLK(clk), .Q(arr[1897]) );
  DFFPOSX1 arr_reg_46__10_ ( .D(n10198), .CLK(clk), .Q(arr[1896]) );
  DFFPOSX1 arr_reg_46__9_ ( .D(n10197), .CLK(clk), .Q(arr[1895]) );
  DFFPOSX1 arr_reg_46__8_ ( .D(n10196), .CLK(clk), .Q(arr[1894]) );
  DFFPOSX1 arr_reg_46__7_ ( .D(n10195), .CLK(clk), .Q(arr[1893]) );
  DFFPOSX1 arr_reg_46__6_ ( .D(n10194), .CLK(clk), .Q(arr[1892]) );
  DFFPOSX1 arr_reg_46__5_ ( .D(n10193), .CLK(clk), .Q(arr[1891]) );
  DFFPOSX1 arr_reg_46__4_ ( .D(n10192), .CLK(clk), .Q(arr[1890]) );
  DFFPOSX1 arr_reg_46__3_ ( .D(n10191), .CLK(clk), .Q(arr[1889]) );
  DFFPOSX1 arr_reg_46__2_ ( .D(n10190), .CLK(clk), .Q(arr[1888]) );
  DFFPOSX1 arr_reg_46__1_ ( .D(n10189), .CLK(clk), .Q(arr[1887]) );
  DFFPOSX1 arr_reg_46__0_ ( .D(n10188), .CLK(clk), .Q(arr[1886]) );
  DFFPOSX1 arr_reg_45__40_ ( .D(n10187), .CLK(clk), .Q(arr[1885]) );
  DFFPOSX1 arr_reg_45__39_ ( .D(n10186), .CLK(clk), .Q(arr[1884]) );
  DFFPOSX1 arr_reg_45__38_ ( .D(n10185), .CLK(clk), .Q(arr[1883]) );
  DFFPOSX1 arr_reg_45__37_ ( .D(n10184), .CLK(clk), .Q(arr[1882]) );
  DFFPOSX1 arr_reg_45__36_ ( .D(n10183), .CLK(clk), .Q(arr[1881]) );
  DFFPOSX1 arr_reg_45__35_ ( .D(n10182), .CLK(clk), .Q(arr[1880]) );
  DFFPOSX1 arr_reg_45__34_ ( .D(n10181), .CLK(clk), .Q(arr[1879]) );
  DFFPOSX1 arr_reg_45__33_ ( .D(n10180), .CLK(clk), .Q(arr[1878]) );
  DFFPOSX1 arr_reg_45__32_ ( .D(n10179), .CLK(clk), .Q(arr[1877]) );
  DFFPOSX1 arr_reg_45__31_ ( .D(n10178), .CLK(clk), .Q(arr[1876]) );
  DFFPOSX1 arr_reg_45__30_ ( .D(n10177), .CLK(clk), .Q(arr[1875]) );
  DFFPOSX1 arr_reg_45__29_ ( .D(n10176), .CLK(clk), .Q(arr[1874]) );
  DFFPOSX1 arr_reg_45__28_ ( .D(n10175), .CLK(clk), .Q(arr[1873]) );
  DFFPOSX1 arr_reg_45__27_ ( .D(n10174), .CLK(clk), .Q(arr[1872]) );
  DFFPOSX1 arr_reg_45__26_ ( .D(n10173), .CLK(clk), .Q(arr[1871]) );
  DFFPOSX1 arr_reg_45__25_ ( .D(n10172), .CLK(clk), .Q(arr[1870]) );
  DFFPOSX1 arr_reg_45__24_ ( .D(n10171), .CLK(clk), .Q(arr[1869]) );
  DFFPOSX1 arr_reg_45__23_ ( .D(n10170), .CLK(clk), .Q(arr[1868]) );
  DFFPOSX1 arr_reg_45__22_ ( .D(n10169), .CLK(clk), .Q(arr[1867]) );
  DFFPOSX1 arr_reg_45__21_ ( .D(n10168), .CLK(clk), .Q(arr[1866]) );
  DFFPOSX1 arr_reg_45__20_ ( .D(n10167), .CLK(clk), .Q(arr[1865]) );
  DFFPOSX1 arr_reg_45__19_ ( .D(n10166), .CLK(clk), .Q(arr[1864]) );
  DFFPOSX1 arr_reg_45__18_ ( .D(n10165), .CLK(clk), .Q(arr[1863]) );
  DFFPOSX1 arr_reg_45__17_ ( .D(n10164), .CLK(clk), .Q(arr[1862]) );
  DFFPOSX1 arr_reg_45__16_ ( .D(n10163), .CLK(clk), .Q(arr[1861]) );
  DFFPOSX1 arr_reg_45__15_ ( .D(n10162), .CLK(clk), .Q(arr[1860]) );
  DFFPOSX1 arr_reg_45__14_ ( .D(n10161), .CLK(clk), .Q(arr[1859]) );
  DFFPOSX1 arr_reg_45__13_ ( .D(n10160), .CLK(clk), .Q(arr[1858]) );
  DFFPOSX1 arr_reg_45__12_ ( .D(n10159), .CLK(clk), .Q(arr[1857]) );
  DFFPOSX1 arr_reg_45__11_ ( .D(n10158), .CLK(clk), .Q(arr[1856]) );
  DFFPOSX1 arr_reg_45__10_ ( .D(n10157), .CLK(clk), .Q(arr[1855]) );
  DFFPOSX1 arr_reg_45__9_ ( .D(n10156), .CLK(clk), .Q(arr[1854]) );
  DFFPOSX1 arr_reg_45__8_ ( .D(n10155), .CLK(clk), .Q(arr[1853]) );
  DFFPOSX1 arr_reg_45__7_ ( .D(n10154), .CLK(clk), .Q(arr[1852]) );
  DFFPOSX1 arr_reg_45__6_ ( .D(n10153), .CLK(clk), .Q(arr[1851]) );
  DFFPOSX1 arr_reg_45__5_ ( .D(n10152), .CLK(clk), .Q(arr[1850]) );
  DFFPOSX1 arr_reg_45__4_ ( .D(n10151), .CLK(clk), .Q(arr[1849]) );
  DFFPOSX1 arr_reg_45__3_ ( .D(n10150), .CLK(clk), .Q(arr[1848]) );
  DFFPOSX1 arr_reg_45__2_ ( .D(n10149), .CLK(clk), .Q(arr[1847]) );
  DFFPOSX1 arr_reg_45__1_ ( .D(n10148), .CLK(clk), .Q(arr[1846]) );
  DFFPOSX1 arr_reg_45__0_ ( .D(n10147), .CLK(clk), .Q(arr[1845]) );
  DFFPOSX1 arr_reg_44__40_ ( .D(n10146), .CLK(clk), .Q(arr[1844]) );
  DFFPOSX1 arr_reg_44__39_ ( .D(n10145), .CLK(clk), .Q(arr[1843]) );
  DFFPOSX1 arr_reg_44__38_ ( .D(n10144), .CLK(clk), .Q(arr[1842]) );
  DFFPOSX1 arr_reg_44__37_ ( .D(n10143), .CLK(clk), .Q(arr[1841]) );
  DFFPOSX1 arr_reg_44__36_ ( .D(n10142), .CLK(clk), .Q(arr[1840]) );
  DFFPOSX1 arr_reg_44__35_ ( .D(n10141), .CLK(clk), .Q(arr[1839]) );
  DFFPOSX1 arr_reg_44__34_ ( .D(n10140), .CLK(clk), .Q(arr[1838]) );
  DFFPOSX1 arr_reg_44__33_ ( .D(n10139), .CLK(clk), .Q(arr[1837]) );
  DFFPOSX1 arr_reg_44__32_ ( .D(n10138), .CLK(clk), .Q(arr[1836]) );
  DFFPOSX1 arr_reg_44__31_ ( .D(n10137), .CLK(clk), .Q(arr[1835]) );
  DFFPOSX1 arr_reg_44__30_ ( .D(n10136), .CLK(clk), .Q(arr[1834]) );
  DFFPOSX1 arr_reg_44__29_ ( .D(n10135), .CLK(clk), .Q(arr[1833]) );
  DFFPOSX1 arr_reg_44__28_ ( .D(n10134), .CLK(clk), .Q(arr[1832]) );
  DFFPOSX1 arr_reg_44__27_ ( .D(n10133), .CLK(clk), .Q(arr[1831]) );
  DFFPOSX1 arr_reg_44__26_ ( .D(n10132), .CLK(clk), .Q(arr[1830]) );
  DFFPOSX1 arr_reg_44__25_ ( .D(n10131), .CLK(clk), .Q(arr[1829]) );
  DFFPOSX1 arr_reg_44__24_ ( .D(n10130), .CLK(clk), .Q(arr[1828]) );
  DFFPOSX1 arr_reg_44__23_ ( .D(n10129), .CLK(clk), .Q(arr[1827]) );
  DFFPOSX1 arr_reg_44__22_ ( .D(n10128), .CLK(clk), .Q(arr[1826]) );
  DFFPOSX1 arr_reg_44__21_ ( .D(n10127), .CLK(clk), .Q(arr[1825]) );
  DFFPOSX1 arr_reg_44__20_ ( .D(n10126), .CLK(clk), .Q(arr[1824]) );
  DFFPOSX1 arr_reg_44__19_ ( .D(n10125), .CLK(clk), .Q(arr[1823]) );
  DFFPOSX1 arr_reg_44__18_ ( .D(n10124), .CLK(clk), .Q(arr[1822]) );
  DFFPOSX1 arr_reg_44__17_ ( .D(n10123), .CLK(clk), .Q(arr[1821]) );
  DFFPOSX1 arr_reg_44__16_ ( .D(n10122), .CLK(clk), .Q(arr[1820]) );
  DFFPOSX1 arr_reg_44__15_ ( .D(n10121), .CLK(clk), .Q(arr[1819]) );
  DFFPOSX1 arr_reg_44__14_ ( .D(n10120), .CLK(clk), .Q(arr[1818]) );
  DFFPOSX1 arr_reg_44__13_ ( .D(n10119), .CLK(clk), .Q(arr[1817]) );
  DFFPOSX1 arr_reg_44__12_ ( .D(n10118), .CLK(clk), .Q(arr[1816]) );
  DFFPOSX1 arr_reg_44__11_ ( .D(n10117), .CLK(clk), .Q(arr[1815]) );
  DFFPOSX1 arr_reg_44__10_ ( .D(n10116), .CLK(clk), .Q(arr[1814]) );
  DFFPOSX1 arr_reg_44__9_ ( .D(n10115), .CLK(clk), .Q(arr[1813]) );
  DFFPOSX1 arr_reg_44__8_ ( .D(n10114), .CLK(clk), .Q(arr[1812]) );
  DFFPOSX1 arr_reg_44__7_ ( .D(n10113), .CLK(clk), .Q(arr[1811]) );
  DFFPOSX1 arr_reg_44__6_ ( .D(n10112), .CLK(clk), .Q(arr[1810]) );
  DFFPOSX1 arr_reg_44__5_ ( .D(n10111), .CLK(clk), .Q(arr[1809]) );
  DFFPOSX1 arr_reg_44__4_ ( .D(n10110), .CLK(clk), .Q(arr[1808]) );
  DFFPOSX1 arr_reg_44__3_ ( .D(n10109), .CLK(clk), .Q(arr[1807]) );
  DFFPOSX1 arr_reg_44__2_ ( .D(n10108), .CLK(clk), .Q(arr[1806]) );
  DFFPOSX1 arr_reg_44__1_ ( .D(n10107), .CLK(clk), .Q(arr[1805]) );
  DFFPOSX1 arr_reg_44__0_ ( .D(n10106), .CLK(clk), .Q(arr[1804]) );
  DFFPOSX1 arr_reg_43__40_ ( .D(n10105), .CLK(clk), .Q(arr[1803]) );
  DFFPOSX1 arr_reg_43__39_ ( .D(n10104), .CLK(clk), .Q(arr[1802]) );
  DFFPOSX1 arr_reg_43__38_ ( .D(n10103), .CLK(clk), .Q(arr[1801]) );
  DFFPOSX1 arr_reg_43__37_ ( .D(n10102), .CLK(clk), .Q(arr[1800]) );
  DFFPOSX1 arr_reg_43__36_ ( .D(n10101), .CLK(clk), .Q(arr[1799]) );
  DFFPOSX1 arr_reg_43__35_ ( .D(n10100), .CLK(clk), .Q(arr[1798]) );
  DFFPOSX1 arr_reg_43__34_ ( .D(n10099), .CLK(clk), .Q(arr[1797]) );
  DFFPOSX1 arr_reg_43__33_ ( .D(n10098), .CLK(clk), .Q(arr[1796]) );
  DFFPOSX1 arr_reg_43__32_ ( .D(n10097), .CLK(clk), .Q(arr[1795]) );
  DFFPOSX1 arr_reg_43__31_ ( .D(n10096), .CLK(clk), .Q(arr[1794]) );
  DFFPOSX1 arr_reg_43__30_ ( .D(n10095), .CLK(clk), .Q(arr[1793]) );
  DFFPOSX1 arr_reg_43__29_ ( .D(n10094), .CLK(clk), .Q(arr[1792]) );
  DFFPOSX1 arr_reg_43__28_ ( .D(n10093), .CLK(clk), .Q(arr[1791]) );
  DFFPOSX1 arr_reg_43__27_ ( .D(n10092), .CLK(clk), .Q(arr[1790]) );
  DFFPOSX1 arr_reg_43__26_ ( .D(n10091), .CLK(clk), .Q(arr[1789]) );
  DFFPOSX1 arr_reg_43__25_ ( .D(n10090), .CLK(clk), .Q(arr[1788]) );
  DFFPOSX1 arr_reg_43__24_ ( .D(n10089), .CLK(clk), .Q(arr[1787]) );
  DFFPOSX1 arr_reg_43__23_ ( .D(n10088), .CLK(clk), .Q(arr[1786]) );
  DFFPOSX1 arr_reg_43__22_ ( .D(n10087), .CLK(clk), .Q(arr[1785]) );
  DFFPOSX1 arr_reg_43__21_ ( .D(n10086), .CLK(clk), .Q(arr[1784]) );
  DFFPOSX1 arr_reg_43__20_ ( .D(n10085), .CLK(clk), .Q(arr[1783]) );
  DFFPOSX1 arr_reg_43__19_ ( .D(n10084), .CLK(clk), .Q(arr[1782]) );
  DFFPOSX1 arr_reg_43__18_ ( .D(n10083), .CLK(clk), .Q(arr[1781]) );
  DFFPOSX1 arr_reg_43__17_ ( .D(n10082), .CLK(clk), .Q(arr[1780]) );
  DFFPOSX1 arr_reg_43__16_ ( .D(n10081), .CLK(clk), .Q(arr[1779]) );
  DFFPOSX1 arr_reg_43__15_ ( .D(n10080), .CLK(clk), .Q(arr[1778]) );
  DFFPOSX1 arr_reg_43__14_ ( .D(n10079), .CLK(clk), .Q(arr[1777]) );
  DFFPOSX1 arr_reg_43__13_ ( .D(n10078), .CLK(clk), .Q(arr[1776]) );
  DFFPOSX1 arr_reg_43__12_ ( .D(n10077), .CLK(clk), .Q(arr[1775]) );
  DFFPOSX1 arr_reg_43__11_ ( .D(n10076), .CLK(clk), .Q(arr[1774]) );
  DFFPOSX1 arr_reg_43__10_ ( .D(n10075), .CLK(clk), .Q(arr[1773]) );
  DFFPOSX1 arr_reg_43__9_ ( .D(n10074), .CLK(clk), .Q(arr[1772]) );
  DFFPOSX1 arr_reg_43__8_ ( .D(n10073), .CLK(clk), .Q(arr[1771]) );
  DFFPOSX1 arr_reg_43__7_ ( .D(n10072), .CLK(clk), .Q(arr[1770]) );
  DFFPOSX1 arr_reg_43__6_ ( .D(n10071), .CLK(clk), .Q(arr[1769]) );
  DFFPOSX1 arr_reg_43__5_ ( .D(n10070), .CLK(clk), .Q(arr[1768]) );
  DFFPOSX1 arr_reg_43__4_ ( .D(n10069), .CLK(clk), .Q(arr[1767]) );
  DFFPOSX1 arr_reg_43__3_ ( .D(n10068), .CLK(clk), .Q(arr[1766]) );
  DFFPOSX1 arr_reg_43__2_ ( .D(n10067), .CLK(clk), .Q(arr[1765]) );
  DFFPOSX1 arr_reg_43__1_ ( .D(n10066), .CLK(clk), .Q(arr[1764]) );
  DFFPOSX1 arr_reg_43__0_ ( .D(n10065), .CLK(clk), .Q(arr[1763]) );
  DFFPOSX1 arr_reg_42__40_ ( .D(n10064), .CLK(clk), .Q(arr[1762]) );
  DFFPOSX1 arr_reg_42__39_ ( .D(n10063), .CLK(clk), .Q(arr[1761]) );
  DFFPOSX1 arr_reg_42__38_ ( .D(n10062), .CLK(clk), .Q(arr[1760]) );
  DFFPOSX1 arr_reg_42__37_ ( .D(n10061), .CLK(clk), .Q(arr[1759]) );
  DFFPOSX1 arr_reg_42__36_ ( .D(n10060), .CLK(clk), .Q(arr[1758]) );
  DFFPOSX1 arr_reg_42__35_ ( .D(n10059), .CLK(clk), .Q(arr[1757]) );
  DFFPOSX1 arr_reg_42__34_ ( .D(n10058), .CLK(clk), .Q(arr[1756]) );
  DFFPOSX1 arr_reg_42__33_ ( .D(n10057), .CLK(clk), .Q(arr[1755]) );
  DFFPOSX1 arr_reg_42__32_ ( .D(n10056), .CLK(clk), .Q(arr[1754]) );
  DFFPOSX1 arr_reg_42__31_ ( .D(n10055), .CLK(clk), .Q(arr[1753]) );
  DFFPOSX1 arr_reg_42__30_ ( .D(n10054), .CLK(clk), .Q(arr[1752]) );
  DFFPOSX1 arr_reg_42__29_ ( .D(n10053), .CLK(clk), .Q(arr[1751]) );
  DFFPOSX1 arr_reg_42__28_ ( .D(n10052), .CLK(clk), .Q(arr[1750]) );
  DFFPOSX1 arr_reg_42__27_ ( .D(n10051), .CLK(clk), .Q(arr[1749]) );
  DFFPOSX1 arr_reg_42__26_ ( .D(n10050), .CLK(clk), .Q(arr[1748]) );
  DFFPOSX1 arr_reg_42__25_ ( .D(n10049), .CLK(clk), .Q(arr[1747]) );
  DFFPOSX1 arr_reg_42__24_ ( .D(n10048), .CLK(clk), .Q(arr[1746]) );
  DFFPOSX1 arr_reg_42__23_ ( .D(n10047), .CLK(clk), .Q(arr[1745]) );
  DFFPOSX1 arr_reg_42__22_ ( .D(n10046), .CLK(clk), .Q(arr[1744]) );
  DFFPOSX1 arr_reg_42__21_ ( .D(n10045), .CLK(clk), .Q(arr[1743]) );
  DFFPOSX1 arr_reg_42__20_ ( .D(n10044), .CLK(clk), .Q(arr[1742]) );
  DFFPOSX1 arr_reg_42__19_ ( .D(n10043), .CLK(clk), .Q(arr[1741]) );
  DFFPOSX1 arr_reg_42__18_ ( .D(n10042), .CLK(clk), .Q(arr[1740]) );
  DFFPOSX1 arr_reg_42__17_ ( .D(n10041), .CLK(clk), .Q(arr[1739]) );
  DFFPOSX1 arr_reg_42__16_ ( .D(n10040), .CLK(clk), .Q(arr[1738]) );
  DFFPOSX1 arr_reg_42__15_ ( .D(n10039), .CLK(clk), .Q(arr[1737]) );
  DFFPOSX1 arr_reg_42__14_ ( .D(n10038), .CLK(clk), .Q(arr[1736]) );
  DFFPOSX1 arr_reg_42__13_ ( .D(n10037), .CLK(clk), .Q(arr[1735]) );
  DFFPOSX1 arr_reg_42__12_ ( .D(n10036), .CLK(clk), .Q(arr[1734]) );
  DFFPOSX1 arr_reg_42__11_ ( .D(n10035), .CLK(clk), .Q(arr[1733]) );
  DFFPOSX1 arr_reg_42__10_ ( .D(n10034), .CLK(clk), .Q(arr[1732]) );
  DFFPOSX1 arr_reg_42__9_ ( .D(n10033), .CLK(clk), .Q(arr[1731]) );
  DFFPOSX1 arr_reg_42__8_ ( .D(n10032), .CLK(clk), .Q(arr[1730]) );
  DFFPOSX1 arr_reg_42__7_ ( .D(n10031), .CLK(clk), .Q(arr[1729]) );
  DFFPOSX1 arr_reg_42__6_ ( .D(n10030), .CLK(clk), .Q(arr[1728]) );
  DFFPOSX1 arr_reg_42__5_ ( .D(n10029), .CLK(clk), .Q(arr[1727]) );
  DFFPOSX1 arr_reg_42__4_ ( .D(n10028), .CLK(clk), .Q(arr[1726]) );
  DFFPOSX1 arr_reg_42__3_ ( .D(n10027), .CLK(clk), .Q(arr[1725]) );
  DFFPOSX1 arr_reg_42__2_ ( .D(n10026), .CLK(clk), .Q(arr[1724]) );
  DFFPOSX1 arr_reg_42__1_ ( .D(n10025), .CLK(clk), .Q(arr[1723]) );
  DFFPOSX1 arr_reg_42__0_ ( .D(n10024), .CLK(clk), .Q(arr[1722]) );
  DFFPOSX1 arr_reg_41__40_ ( .D(n10023), .CLK(clk), .Q(arr[1721]) );
  DFFPOSX1 arr_reg_41__39_ ( .D(n10022), .CLK(clk), .Q(arr[1720]) );
  DFFPOSX1 arr_reg_41__38_ ( .D(n10021), .CLK(clk), .Q(arr[1719]) );
  DFFPOSX1 arr_reg_41__37_ ( .D(n10020), .CLK(clk), .Q(arr[1718]) );
  DFFPOSX1 arr_reg_41__36_ ( .D(n10019), .CLK(clk), .Q(arr[1717]) );
  DFFPOSX1 arr_reg_41__35_ ( .D(n10018), .CLK(clk), .Q(arr[1716]) );
  DFFPOSX1 arr_reg_41__34_ ( .D(n10017), .CLK(clk), .Q(arr[1715]) );
  DFFPOSX1 arr_reg_41__33_ ( .D(n10016), .CLK(clk), .Q(arr[1714]) );
  DFFPOSX1 arr_reg_41__32_ ( .D(n10015), .CLK(clk), .Q(arr[1713]) );
  DFFPOSX1 arr_reg_41__31_ ( .D(n10014), .CLK(clk), .Q(arr[1712]) );
  DFFPOSX1 arr_reg_41__30_ ( .D(n10013), .CLK(clk), .Q(arr[1711]) );
  DFFPOSX1 arr_reg_41__29_ ( .D(n10012), .CLK(clk), .Q(arr[1710]) );
  DFFPOSX1 arr_reg_41__28_ ( .D(n10011), .CLK(clk), .Q(arr[1709]) );
  DFFPOSX1 arr_reg_41__27_ ( .D(n10010), .CLK(clk), .Q(arr[1708]) );
  DFFPOSX1 arr_reg_41__26_ ( .D(n10009), .CLK(clk), .Q(arr[1707]) );
  DFFPOSX1 arr_reg_41__25_ ( .D(n10008), .CLK(clk), .Q(arr[1706]) );
  DFFPOSX1 arr_reg_41__24_ ( .D(n10007), .CLK(clk), .Q(arr[1705]) );
  DFFPOSX1 arr_reg_41__23_ ( .D(n10006), .CLK(clk), .Q(arr[1704]) );
  DFFPOSX1 arr_reg_41__22_ ( .D(n10005), .CLK(clk), .Q(arr[1703]) );
  DFFPOSX1 arr_reg_41__21_ ( .D(n10004), .CLK(clk), .Q(arr[1702]) );
  DFFPOSX1 arr_reg_41__20_ ( .D(n10003), .CLK(clk), .Q(arr[1701]) );
  DFFPOSX1 arr_reg_41__19_ ( .D(n10002), .CLK(clk), .Q(arr[1700]) );
  DFFPOSX1 arr_reg_41__18_ ( .D(n10001), .CLK(clk), .Q(arr[1699]) );
  DFFPOSX1 arr_reg_41__17_ ( .D(n10000), .CLK(clk), .Q(arr[1698]) );
  DFFPOSX1 arr_reg_41__16_ ( .D(n9999), .CLK(clk), .Q(arr[1697]) );
  DFFPOSX1 arr_reg_41__15_ ( .D(n9998), .CLK(clk), .Q(arr[1696]) );
  DFFPOSX1 arr_reg_41__14_ ( .D(n9997), .CLK(clk), .Q(arr[1695]) );
  DFFPOSX1 arr_reg_41__13_ ( .D(n9996), .CLK(clk), .Q(arr[1694]) );
  DFFPOSX1 arr_reg_41__12_ ( .D(n9995), .CLK(clk), .Q(arr[1693]) );
  DFFPOSX1 arr_reg_41__11_ ( .D(n9994), .CLK(clk), .Q(arr[1692]) );
  DFFPOSX1 arr_reg_41__10_ ( .D(n9993), .CLK(clk), .Q(arr[1691]) );
  DFFPOSX1 arr_reg_41__9_ ( .D(n9992), .CLK(clk), .Q(arr[1690]) );
  DFFPOSX1 arr_reg_41__8_ ( .D(n9991), .CLK(clk), .Q(arr[1689]) );
  DFFPOSX1 arr_reg_41__7_ ( .D(n9990), .CLK(clk), .Q(arr[1688]) );
  DFFPOSX1 arr_reg_41__6_ ( .D(n9989), .CLK(clk), .Q(arr[1687]) );
  DFFPOSX1 arr_reg_41__5_ ( .D(n9988), .CLK(clk), .Q(arr[1686]) );
  DFFPOSX1 arr_reg_41__4_ ( .D(n9987), .CLK(clk), .Q(arr[1685]) );
  DFFPOSX1 arr_reg_41__3_ ( .D(n9986), .CLK(clk), .Q(arr[1684]) );
  DFFPOSX1 arr_reg_41__2_ ( .D(n9985), .CLK(clk), .Q(arr[1683]) );
  DFFPOSX1 arr_reg_41__1_ ( .D(n9984), .CLK(clk), .Q(arr[1682]) );
  DFFPOSX1 arr_reg_41__0_ ( .D(n9983), .CLK(clk), .Q(arr[1681]) );
  DFFPOSX1 arr_reg_40__40_ ( .D(n9982), .CLK(clk), .Q(arr[1680]) );
  DFFPOSX1 arr_reg_40__39_ ( .D(n9981), .CLK(clk), .Q(arr[1679]) );
  DFFPOSX1 arr_reg_40__38_ ( .D(n9980), .CLK(clk), .Q(arr[1678]) );
  DFFPOSX1 arr_reg_40__37_ ( .D(n9979), .CLK(clk), .Q(arr[1677]) );
  DFFPOSX1 arr_reg_40__36_ ( .D(n9978), .CLK(clk), .Q(arr[1676]) );
  DFFPOSX1 arr_reg_40__35_ ( .D(n9977), .CLK(clk), .Q(arr[1675]) );
  DFFPOSX1 arr_reg_40__34_ ( .D(n9976), .CLK(clk), .Q(arr[1674]) );
  DFFPOSX1 arr_reg_40__33_ ( .D(n9975), .CLK(clk), .Q(arr[1673]) );
  DFFPOSX1 arr_reg_40__32_ ( .D(n9974), .CLK(clk), .Q(arr[1672]) );
  DFFPOSX1 arr_reg_40__31_ ( .D(n9973), .CLK(clk), .Q(arr[1671]) );
  DFFPOSX1 arr_reg_40__30_ ( .D(n9972), .CLK(clk), .Q(arr[1670]) );
  DFFPOSX1 arr_reg_40__29_ ( .D(n9971), .CLK(clk), .Q(arr[1669]) );
  DFFPOSX1 arr_reg_40__28_ ( .D(n9970), .CLK(clk), .Q(arr[1668]) );
  DFFPOSX1 arr_reg_40__27_ ( .D(n9969), .CLK(clk), .Q(arr[1667]) );
  DFFPOSX1 arr_reg_40__26_ ( .D(n9968), .CLK(clk), .Q(arr[1666]) );
  DFFPOSX1 arr_reg_40__25_ ( .D(n9967), .CLK(clk), .Q(arr[1665]) );
  DFFPOSX1 arr_reg_40__24_ ( .D(n9966), .CLK(clk), .Q(arr[1664]) );
  DFFPOSX1 arr_reg_40__23_ ( .D(n9965), .CLK(clk), .Q(arr[1663]) );
  DFFPOSX1 arr_reg_40__22_ ( .D(n9964), .CLK(clk), .Q(arr[1662]) );
  DFFPOSX1 arr_reg_40__21_ ( .D(n9963), .CLK(clk), .Q(arr[1661]) );
  DFFPOSX1 arr_reg_40__20_ ( .D(n9962), .CLK(clk), .Q(arr[1660]) );
  DFFPOSX1 arr_reg_40__19_ ( .D(n9961), .CLK(clk), .Q(arr[1659]) );
  DFFPOSX1 arr_reg_40__18_ ( .D(n9960), .CLK(clk), .Q(arr[1658]) );
  DFFPOSX1 arr_reg_40__17_ ( .D(n9959), .CLK(clk), .Q(arr[1657]) );
  DFFPOSX1 arr_reg_40__16_ ( .D(n9958), .CLK(clk), .Q(arr[1656]) );
  DFFPOSX1 arr_reg_40__15_ ( .D(n9957), .CLK(clk), .Q(arr[1655]) );
  DFFPOSX1 arr_reg_40__14_ ( .D(n9956), .CLK(clk), .Q(arr[1654]) );
  DFFPOSX1 arr_reg_40__13_ ( .D(n9955), .CLK(clk), .Q(arr[1653]) );
  DFFPOSX1 arr_reg_40__12_ ( .D(n9954), .CLK(clk), .Q(arr[1652]) );
  DFFPOSX1 arr_reg_40__11_ ( .D(n9953), .CLK(clk), .Q(arr[1651]) );
  DFFPOSX1 arr_reg_40__10_ ( .D(n9952), .CLK(clk), .Q(arr[1650]) );
  DFFPOSX1 arr_reg_40__9_ ( .D(n9951), .CLK(clk), .Q(arr[1649]) );
  DFFPOSX1 arr_reg_40__8_ ( .D(n9950), .CLK(clk), .Q(arr[1648]) );
  DFFPOSX1 arr_reg_40__7_ ( .D(n9949), .CLK(clk), .Q(arr[1647]) );
  DFFPOSX1 arr_reg_40__6_ ( .D(n9948), .CLK(clk), .Q(arr[1646]) );
  DFFPOSX1 arr_reg_40__5_ ( .D(n9947), .CLK(clk), .Q(arr[1645]) );
  DFFPOSX1 arr_reg_40__4_ ( .D(n9946), .CLK(clk), .Q(arr[1644]) );
  DFFPOSX1 arr_reg_40__3_ ( .D(n9945), .CLK(clk), .Q(arr[1643]) );
  DFFPOSX1 arr_reg_40__2_ ( .D(n9944), .CLK(clk), .Q(arr[1642]) );
  DFFPOSX1 arr_reg_40__1_ ( .D(n9943), .CLK(clk), .Q(arr[1641]) );
  DFFPOSX1 arr_reg_40__0_ ( .D(n9942), .CLK(clk), .Q(arr[1640]) );
  DFFPOSX1 arr_reg_39__40_ ( .D(n9941), .CLK(clk), .Q(arr[1639]) );
  DFFPOSX1 arr_reg_39__39_ ( .D(n9940), .CLK(clk), .Q(arr[1638]) );
  DFFPOSX1 arr_reg_39__38_ ( .D(n9939), .CLK(clk), .Q(arr[1637]) );
  DFFPOSX1 arr_reg_39__37_ ( .D(n9938), .CLK(clk), .Q(arr[1636]) );
  DFFPOSX1 arr_reg_39__36_ ( .D(n9937), .CLK(clk), .Q(arr[1635]) );
  DFFPOSX1 arr_reg_39__35_ ( .D(n9936), .CLK(clk), .Q(arr[1634]) );
  DFFPOSX1 arr_reg_39__34_ ( .D(n9935), .CLK(clk), .Q(arr[1633]) );
  DFFPOSX1 arr_reg_39__33_ ( .D(n9934), .CLK(clk), .Q(arr[1632]) );
  DFFPOSX1 arr_reg_39__32_ ( .D(n9933), .CLK(clk), .Q(arr[1631]) );
  DFFPOSX1 arr_reg_39__31_ ( .D(n9932), .CLK(clk), .Q(arr[1630]) );
  DFFPOSX1 arr_reg_39__30_ ( .D(n9931), .CLK(clk), .Q(arr[1629]) );
  DFFPOSX1 arr_reg_39__29_ ( .D(n9930), .CLK(clk), .Q(arr[1628]) );
  DFFPOSX1 arr_reg_39__28_ ( .D(n9929), .CLK(clk), .Q(arr[1627]) );
  DFFPOSX1 arr_reg_39__27_ ( .D(n9928), .CLK(clk), .Q(arr[1626]) );
  DFFPOSX1 arr_reg_39__26_ ( .D(n9927), .CLK(clk), .Q(arr[1625]) );
  DFFPOSX1 arr_reg_39__25_ ( .D(n9926), .CLK(clk), .Q(arr[1624]) );
  DFFPOSX1 arr_reg_39__24_ ( .D(n9925), .CLK(clk), .Q(arr[1623]) );
  DFFPOSX1 arr_reg_39__23_ ( .D(n9924), .CLK(clk), .Q(arr[1622]) );
  DFFPOSX1 arr_reg_39__22_ ( .D(n9923), .CLK(clk), .Q(arr[1621]) );
  DFFPOSX1 arr_reg_39__21_ ( .D(n9922), .CLK(clk), .Q(arr[1620]) );
  DFFPOSX1 arr_reg_39__20_ ( .D(n9921), .CLK(clk), .Q(arr[1619]) );
  DFFPOSX1 arr_reg_39__19_ ( .D(n9920), .CLK(clk), .Q(arr[1618]) );
  DFFPOSX1 arr_reg_39__18_ ( .D(n9919), .CLK(clk), .Q(arr[1617]) );
  DFFPOSX1 arr_reg_39__17_ ( .D(n9918), .CLK(clk), .Q(arr[1616]) );
  DFFPOSX1 arr_reg_39__16_ ( .D(n9917), .CLK(clk), .Q(arr[1615]) );
  DFFPOSX1 arr_reg_39__15_ ( .D(n9916), .CLK(clk), .Q(arr[1614]) );
  DFFPOSX1 arr_reg_39__14_ ( .D(n9915), .CLK(clk), .Q(arr[1613]) );
  DFFPOSX1 arr_reg_39__13_ ( .D(n9914), .CLK(clk), .Q(arr[1612]) );
  DFFPOSX1 arr_reg_39__12_ ( .D(n9913), .CLK(clk), .Q(arr[1611]) );
  DFFPOSX1 arr_reg_39__11_ ( .D(n9912), .CLK(clk), .Q(arr[1610]) );
  DFFPOSX1 arr_reg_39__10_ ( .D(n9911), .CLK(clk), .Q(arr[1609]) );
  DFFPOSX1 arr_reg_39__9_ ( .D(n9910), .CLK(clk), .Q(arr[1608]) );
  DFFPOSX1 arr_reg_39__8_ ( .D(n9909), .CLK(clk), .Q(arr[1607]) );
  DFFPOSX1 arr_reg_39__7_ ( .D(n9908), .CLK(clk), .Q(arr[1606]) );
  DFFPOSX1 arr_reg_39__6_ ( .D(n9907), .CLK(clk), .Q(arr[1605]) );
  DFFPOSX1 arr_reg_39__5_ ( .D(n9906), .CLK(clk), .Q(arr[1604]) );
  DFFPOSX1 arr_reg_39__4_ ( .D(n9905), .CLK(clk), .Q(arr[1603]) );
  DFFPOSX1 arr_reg_39__3_ ( .D(n9904), .CLK(clk), .Q(arr[1602]) );
  DFFPOSX1 arr_reg_39__2_ ( .D(n9903), .CLK(clk), .Q(arr[1601]) );
  DFFPOSX1 arr_reg_39__1_ ( .D(n9902), .CLK(clk), .Q(arr[1600]) );
  DFFPOSX1 arr_reg_39__0_ ( .D(n9901), .CLK(clk), .Q(arr[1599]) );
  DFFPOSX1 arr_reg_38__40_ ( .D(n9900), .CLK(clk), .Q(arr[1598]) );
  DFFPOSX1 arr_reg_38__39_ ( .D(n9899), .CLK(clk), .Q(arr[1597]) );
  DFFPOSX1 arr_reg_38__38_ ( .D(n9898), .CLK(clk), .Q(arr[1596]) );
  DFFPOSX1 arr_reg_38__37_ ( .D(n9897), .CLK(clk), .Q(arr[1595]) );
  DFFPOSX1 arr_reg_38__36_ ( .D(n9896), .CLK(clk), .Q(arr[1594]) );
  DFFPOSX1 arr_reg_38__35_ ( .D(n9895), .CLK(clk), .Q(arr[1593]) );
  DFFPOSX1 arr_reg_38__34_ ( .D(n9894), .CLK(clk), .Q(arr[1592]) );
  DFFPOSX1 arr_reg_38__33_ ( .D(n9893), .CLK(clk), .Q(arr[1591]) );
  DFFPOSX1 arr_reg_38__32_ ( .D(n9892), .CLK(clk), .Q(arr[1590]) );
  DFFPOSX1 arr_reg_38__31_ ( .D(n9891), .CLK(clk), .Q(arr[1589]) );
  DFFPOSX1 arr_reg_38__30_ ( .D(n9890), .CLK(clk), .Q(arr[1588]) );
  DFFPOSX1 arr_reg_38__29_ ( .D(n9889), .CLK(clk), .Q(arr[1587]) );
  DFFPOSX1 arr_reg_38__28_ ( .D(n9888), .CLK(clk), .Q(arr[1586]) );
  DFFPOSX1 arr_reg_38__27_ ( .D(n9887), .CLK(clk), .Q(arr[1585]) );
  DFFPOSX1 arr_reg_38__26_ ( .D(n9886), .CLK(clk), .Q(arr[1584]) );
  DFFPOSX1 arr_reg_38__25_ ( .D(n9885), .CLK(clk), .Q(arr[1583]) );
  DFFPOSX1 arr_reg_38__24_ ( .D(n9884), .CLK(clk), .Q(arr[1582]) );
  DFFPOSX1 arr_reg_38__23_ ( .D(n9883), .CLK(clk), .Q(arr[1581]) );
  DFFPOSX1 arr_reg_38__22_ ( .D(n9882), .CLK(clk), .Q(arr[1580]) );
  DFFPOSX1 arr_reg_38__21_ ( .D(n9881), .CLK(clk), .Q(arr[1579]) );
  DFFPOSX1 arr_reg_38__20_ ( .D(n9880), .CLK(clk), .Q(arr[1578]) );
  DFFPOSX1 arr_reg_38__19_ ( .D(n9879), .CLK(clk), .Q(arr[1577]) );
  DFFPOSX1 arr_reg_38__18_ ( .D(n9878), .CLK(clk), .Q(arr[1576]) );
  DFFPOSX1 arr_reg_38__17_ ( .D(n9877), .CLK(clk), .Q(arr[1575]) );
  DFFPOSX1 arr_reg_38__16_ ( .D(n9876), .CLK(clk), .Q(arr[1574]) );
  DFFPOSX1 arr_reg_38__15_ ( .D(n9875), .CLK(clk), .Q(arr[1573]) );
  DFFPOSX1 arr_reg_38__14_ ( .D(n9874), .CLK(clk), .Q(arr[1572]) );
  DFFPOSX1 arr_reg_38__13_ ( .D(n9873), .CLK(clk), .Q(arr[1571]) );
  DFFPOSX1 arr_reg_38__12_ ( .D(n9872), .CLK(clk), .Q(arr[1570]) );
  DFFPOSX1 arr_reg_38__11_ ( .D(n9871), .CLK(clk), .Q(arr[1569]) );
  DFFPOSX1 arr_reg_38__10_ ( .D(n9870), .CLK(clk), .Q(arr[1568]) );
  DFFPOSX1 arr_reg_38__9_ ( .D(n9869), .CLK(clk), .Q(arr[1567]) );
  DFFPOSX1 arr_reg_38__8_ ( .D(n9868), .CLK(clk), .Q(arr[1566]) );
  DFFPOSX1 arr_reg_38__7_ ( .D(n9867), .CLK(clk), .Q(arr[1565]) );
  DFFPOSX1 arr_reg_38__6_ ( .D(n9866), .CLK(clk), .Q(arr[1564]) );
  DFFPOSX1 arr_reg_38__5_ ( .D(n9865), .CLK(clk), .Q(arr[1563]) );
  DFFPOSX1 arr_reg_38__4_ ( .D(n9864), .CLK(clk), .Q(arr[1562]) );
  DFFPOSX1 arr_reg_38__3_ ( .D(n9863), .CLK(clk), .Q(arr[1561]) );
  DFFPOSX1 arr_reg_38__2_ ( .D(n9862), .CLK(clk), .Q(arr[1560]) );
  DFFPOSX1 arr_reg_38__1_ ( .D(n9861), .CLK(clk), .Q(arr[1559]) );
  DFFPOSX1 arr_reg_38__0_ ( .D(n9860), .CLK(clk), .Q(arr[1558]) );
  DFFPOSX1 arr_reg_37__40_ ( .D(n9859), .CLK(clk), .Q(arr[1557]) );
  DFFPOSX1 arr_reg_37__39_ ( .D(n9858), .CLK(clk), .Q(arr[1556]) );
  DFFPOSX1 arr_reg_37__38_ ( .D(n9857), .CLK(clk), .Q(arr[1555]) );
  DFFPOSX1 arr_reg_37__37_ ( .D(n9856), .CLK(clk), .Q(arr[1554]) );
  DFFPOSX1 arr_reg_37__36_ ( .D(n9855), .CLK(clk), .Q(arr[1553]) );
  DFFPOSX1 arr_reg_37__35_ ( .D(n9854), .CLK(clk), .Q(arr[1552]) );
  DFFPOSX1 arr_reg_37__34_ ( .D(n9853), .CLK(clk), .Q(arr[1551]) );
  DFFPOSX1 arr_reg_37__33_ ( .D(n9852), .CLK(clk), .Q(arr[1550]) );
  DFFPOSX1 arr_reg_37__32_ ( .D(n9851), .CLK(clk), .Q(arr[1549]) );
  DFFPOSX1 arr_reg_37__31_ ( .D(n9850), .CLK(clk), .Q(arr[1548]) );
  DFFPOSX1 arr_reg_37__30_ ( .D(n9849), .CLK(clk), .Q(arr[1547]) );
  DFFPOSX1 arr_reg_37__29_ ( .D(n9848), .CLK(clk), .Q(arr[1546]) );
  DFFPOSX1 arr_reg_37__28_ ( .D(n9847), .CLK(clk), .Q(arr[1545]) );
  DFFPOSX1 arr_reg_37__27_ ( .D(n9846), .CLK(clk), .Q(arr[1544]) );
  DFFPOSX1 arr_reg_37__26_ ( .D(n9845), .CLK(clk), .Q(arr[1543]) );
  DFFPOSX1 arr_reg_37__25_ ( .D(n9844), .CLK(clk), .Q(arr[1542]) );
  DFFPOSX1 arr_reg_37__24_ ( .D(n9843), .CLK(clk), .Q(arr[1541]) );
  DFFPOSX1 arr_reg_37__23_ ( .D(n9842), .CLK(clk), .Q(arr[1540]) );
  DFFPOSX1 arr_reg_37__22_ ( .D(n9841), .CLK(clk), .Q(arr[1539]) );
  DFFPOSX1 arr_reg_37__21_ ( .D(n9840), .CLK(clk), .Q(arr[1538]) );
  DFFPOSX1 arr_reg_37__20_ ( .D(n9839), .CLK(clk), .Q(arr[1537]) );
  DFFPOSX1 arr_reg_37__19_ ( .D(n9838), .CLK(clk), .Q(arr[1536]) );
  DFFPOSX1 arr_reg_37__18_ ( .D(n9837), .CLK(clk), .Q(arr[1535]) );
  DFFPOSX1 arr_reg_37__17_ ( .D(n9836), .CLK(clk), .Q(arr[1534]) );
  DFFPOSX1 arr_reg_37__16_ ( .D(n9835), .CLK(clk), .Q(arr[1533]) );
  DFFPOSX1 arr_reg_37__15_ ( .D(n9834), .CLK(clk), .Q(arr[1532]) );
  DFFPOSX1 arr_reg_37__14_ ( .D(n9833), .CLK(clk), .Q(arr[1531]) );
  DFFPOSX1 arr_reg_37__13_ ( .D(n9832), .CLK(clk), .Q(arr[1530]) );
  DFFPOSX1 arr_reg_37__12_ ( .D(n9831), .CLK(clk), .Q(arr[1529]) );
  DFFPOSX1 arr_reg_37__11_ ( .D(n9830), .CLK(clk), .Q(arr[1528]) );
  DFFPOSX1 arr_reg_37__10_ ( .D(n9829), .CLK(clk), .Q(arr[1527]) );
  DFFPOSX1 arr_reg_37__9_ ( .D(n9828), .CLK(clk), .Q(arr[1526]) );
  DFFPOSX1 arr_reg_37__8_ ( .D(n9827), .CLK(clk), .Q(arr[1525]) );
  DFFPOSX1 arr_reg_37__7_ ( .D(n9826), .CLK(clk), .Q(arr[1524]) );
  DFFPOSX1 arr_reg_37__6_ ( .D(n9825), .CLK(clk), .Q(arr[1523]) );
  DFFPOSX1 arr_reg_37__5_ ( .D(n9824), .CLK(clk), .Q(arr[1522]) );
  DFFPOSX1 arr_reg_37__4_ ( .D(n9823), .CLK(clk), .Q(arr[1521]) );
  DFFPOSX1 arr_reg_37__3_ ( .D(n9822), .CLK(clk), .Q(arr[1520]) );
  DFFPOSX1 arr_reg_37__2_ ( .D(n9821), .CLK(clk), .Q(arr[1519]) );
  DFFPOSX1 arr_reg_37__1_ ( .D(n9820), .CLK(clk), .Q(arr[1518]) );
  DFFPOSX1 arr_reg_37__0_ ( .D(n9819), .CLK(clk), .Q(arr[1517]) );
  DFFPOSX1 arr_reg_36__40_ ( .D(n9818), .CLK(clk), .Q(arr[1516]) );
  DFFPOSX1 arr_reg_36__39_ ( .D(n9817), .CLK(clk), .Q(arr[1515]) );
  DFFPOSX1 arr_reg_36__38_ ( .D(n9816), .CLK(clk), .Q(arr[1514]) );
  DFFPOSX1 arr_reg_36__37_ ( .D(n9815), .CLK(clk), .Q(arr[1513]) );
  DFFPOSX1 arr_reg_36__36_ ( .D(n9814), .CLK(clk), .Q(arr[1512]) );
  DFFPOSX1 arr_reg_36__35_ ( .D(n9813), .CLK(clk), .Q(arr[1511]) );
  DFFPOSX1 arr_reg_36__34_ ( .D(n9812), .CLK(clk), .Q(arr[1510]) );
  DFFPOSX1 arr_reg_36__33_ ( .D(n9811), .CLK(clk), .Q(arr[1509]) );
  DFFPOSX1 arr_reg_36__32_ ( .D(n9810), .CLK(clk), .Q(arr[1508]) );
  DFFPOSX1 arr_reg_36__31_ ( .D(n9809), .CLK(clk), .Q(arr[1507]) );
  DFFPOSX1 arr_reg_36__30_ ( .D(n9808), .CLK(clk), .Q(arr[1506]) );
  DFFPOSX1 arr_reg_36__29_ ( .D(n9807), .CLK(clk), .Q(arr[1505]) );
  DFFPOSX1 arr_reg_36__28_ ( .D(n9806), .CLK(clk), .Q(arr[1504]) );
  DFFPOSX1 arr_reg_36__27_ ( .D(n9805), .CLK(clk), .Q(arr[1503]) );
  DFFPOSX1 arr_reg_36__26_ ( .D(n9804), .CLK(clk), .Q(arr[1502]) );
  DFFPOSX1 arr_reg_36__25_ ( .D(n9803), .CLK(clk), .Q(arr[1501]) );
  DFFPOSX1 arr_reg_36__24_ ( .D(n9802), .CLK(clk), .Q(arr[1500]) );
  DFFPOSX1 arr_reg_36__23_ ( .D(n9801), .CLK(clk), .Q(arr[1499]) );
  DFFPOSX1 arr_reg_36__22_ ( .D(n9800), .CLK(clk), .Q(arr[1498]) );
  DFFPOSX1 arr_reg_36__21_ ( .D(n9799), .CLK(clk), .Q(arr[1497]) );
  DFFPOSX1 arr_reg_36__20_ ( .D(n9798), .CLK(clk), .Q(arr[1496]) );
  DFFPOSX1 arr_reg_36__19_ ( .D(n9797), .CLK(clk), .Q(arr[1495]) );
  DFFPOSX1 arr_reg_36__18_ ( .D(n9796), .CLK(clk), .Q(arr[1494]) );
  DFFPOSX1 arr_reg_36__17_ ( .D(n9795), .CLK(clk), .Q(arr[1493]) );
  DFFPOSX1 arr_reg_36__16_ ( .D(n9794), .CLK(clk), .Q(arr[1492]) );
  DFFPOSX1 arr_reg_36__15_ ( .D(n9793), .CLK(clk), .Q(arr[1491]) );
  DFFPOSX1 arr_reg_36__14_ ( .D(n9792), .CLK(clk), .Q(arr[1490]) );
  DFFPOSX1 arr_reg_36__13_ ( .D(n9791), .CLK(clk), .Q(arr[1489]) );
  DFFPOSX1 arr_reg_36__12_ ( .D(n9790), .CLK(clk), .Q(arr[1488]) );
  DFFPOSX1 arr_reg_36__11_ ( .D(n9789), .CLK(clk), .Q(arr[1487]) );
  DFFPOSX1 arr_reg_36__10_ ( .D(n9788), .CLK(clk), .Q(arr[1486]) );
  DFFPOSX1 arr_reg_36__9_ ( .D(n9787), .CLK(clk), .Q(arr[1485]) );
  DFFPOSX1 arr_reg_36__8_ ( .D(n9786), .CLK(clk), .Q(arr[1484]) );
  DFFPOSX1 arr_reg_36__7_ ( .D(n9785), .CLK(clk), .Q(arr[1483]) );
  DFFPOSX1 arr_reg_36__6_ ( .D(n9784), .CLK(clk), .Q(arr[1482]) );
  DFFPOSX1 arr_reg_36__5_ ( .D(n9783), .CLK(clk), .Q(arr[1481]) );
  DFFPOSX1 arr_reg_36__4_ ( .D(n9782), .CLK(clk), .Q(arr[1480]) );
  DFFPOSX1 arr_reg_36__3_ ( .D(n9781), .CLK(clk), .Q(arr[1479]) );
  DFFPOSX1 arr_reg_36__2_ ( .D(n9780), .CLK(clk), .Q(arr[1478]) );
  DFFPOSX1 arr_reg_36__1_ ( .D(n9779), .CLK(clk), .Q(arr[1477]) );
  DFFPOSX1 arr_reg_36__0_ ( .D(n9778), .CLK(clk), .Q(arr[1476]) );
  DFFPOSX1 arr_reg_35__40_ ( .D(n9777), .CLK(clk), .Q(arr[1475]) );
  DFFPOSX1 arr_reg_35__39_ ( .D(n9776), .CLK(clk), .Q(arr[1474]) );
  DFFPOSX1 arr_reg_35__38_ ( .D(n9775), .CLK(clk), .Q(arr[1473]) );
  DFFPOSX1 arr_reg_35__37_ ( .D(n9774), .CLK(clk), .Q(arr[1472]) );
  DFFPOSX1 arr_reg_35__36_ ( .D(n9773), .CLK(clk), .Q(arr[1471]) );
  DFFPOSX1 arr_reg_35__35_ ( .D(n9772), .CLK(clk), .Q(arr[1470]) );
  DFFPOSX1 arr_reg_35__34_ ( .D(n9771), .CLK(clk), .Q(arr[1469]) );
  DFFPOSX1 arr_reg_35__33_ ( .D(n9770), .CLK(clk), .Q(arr[1468]) );
  DFFPOSX1 arr_reg_35__32_ ( .D(n9769), .CLK(clk), .Q(arr[1467]) );
  DFFPOSX1 arr_reg_35__31_ ( .D(n9768), .CLK(clk), .Q(arr[1466]) );
  DFFPOSX1 arr_reg_35__30_ ( .D(n9767), .CLK(clk), .Q(arr[1465]) );
  DFFPOSX1 arr_reg_35__29_ ( .D(n9766), .CLK(clk), .Q(arr[1464]) );
  DFFPOSX1 arr_reg_35__28_ ( .D(n9765), .CLK(clk), .Q(arr[1463]) );
  DFFPOSX1 arr_reg_35__27_ ( .D(n9764), .CLK(clk), .Q(arr[1462]) );
  DFFPOSX1 arr_reg_35__26_ ( .D(n9763), .CLK(clk), .Q(arr[1461]) );
  DFFPOSX1 arr_reg_35__25_ ( .D(n9762), .CLK(clk), .Q(arr[1460]) );
  DFFPOSX1 arr_reg_35__24_ ( .D(n9761), .CLK(clk), .Q(arr[1459]) );
  DFFPOSX1 arr_reg_35__23_ ( .D(n9760), .CLK(clk), .Q(arr[1458]) );
  DFFPOSX1 arr_reg_35__22_ ( .D(n9759), .CLK(clk), .Q(arr[1457]) );
  DFFPOSX1 arr_reg_35__21_ ( .D(n9758), .CLK(clk), .Q(arr[1456]) );
  DFFPOSX1 arr_reg_35__20_ ( .D(n9757), .CLK(clk), .Q(arr[1455]) );
  DFFPOSX1 arr_reg_35__19_ ( .D(n9756), .CLK(clk), .Q(arr[1454]) );
  DFFPOSX1 arr_reg_35__18_ ( .D(n9755), .CLK(clk), .Q(arr[1453]) );
  DFFPOSX1 arr_reg_35__17_ ( .D(n9754), .CLK(clk), .Q(arr[1452]) );
  DFFPOSX1 arr_reg_35__16_ ( .D(n9753), .CLK(clk), .Q(arr[1451]) );
  DFFPOSX1 arr_reg_35__15_ ( .D(n9752), .CLK(clk), .Q(arr[1450]) );
  DFFPOSX1 arr_reg_35__14_ ( .D(n9751), .CLK(clk), .Q(arr[1449]) );
  DFFPOSX1 arr_reg_35__13_ ( .D(n9750), .CLK(clk), .Q(arr[1448]) );
  DFFPOSX1 arr_reg_35__12_ ( .D(n9749), .CLK(clk), .Q(arr[1447]) );
  DFFPOSX1 arr_reg_35__11_ ( .D(n9748), .CLK(clk), .Q(arr[1446]) );
  DFFPOSX1 arr_reg_35__10_ ( .D(n9747), .CLK(clk), .Q(arr[1445]) );
  DFFPOSX1 arr_reg_35__9_ ( .D(n9746), .CLK(clk), .Q(arr[1444]) );
  DFFPOSX1 arr_reg_35__8_ ( .D(n9745), .CLK(clk), .Q(arr[1443]) );
  DFFPOSX1 arr_reg_35__7_ ( .D(n9744), .CLK(clk), .Q(arr[1442]) );
  DFFPOSX1 arr_reg_35__6_ ( .D(n9743), .CLK(clk), .Q(arr[1441]) );
  DFFPOSX1 arr_reg_35__5_ ( .D(n9742), .CLK(clk), .Q(arr[1440]) );
  DFFPOSX1 arr_reg_35__4_ ( .D(n9741), .CLK(clk), .Q(arr[1439]) );
  DFFPOSX1 arr_reg_35__3_ ( .D(n9740), .CLK(clk), .Q(arr[1438]) );
  DFFPOSX1 arr_reg_35__2_ ( .D(n9739), .CLK(clk), .Q(arr[1437]) );
  DFFPOSX1 arr_reg_35__1_ ( .D(n9738), .CLK(clk), .Q(arr[1436]) );
  DFFPOSX1 arr_reg_35__0_ ( .D(n9737), .CLK(clk), .Q(arr[1435]) );
  DFFPOSX1 arr_reg_34__40_ ( .D(n9736), .CLK(clk), .Q(arr[1434]) );
  DFFPOSX1 arr_reg_34__39_ ( .D(n9735), .CLK(clk), .Q(arr[1433]) );
  DFFPOSX1 arr_reg_34__38_ ( .D(n9734), .CLK(clk), .Q(arr[1432]) );
  DFFPOSX1 arr_reg_34__37_ ( .D(n9733), .CLK(clk), .Q(arr[1431]) );
  DFFPOSX1 arr_reg_34__36_ ( .D(n9732), .CLK(clk), .Q(arr[1430]) );
  DFFPOSX1 arr_reg_34__35_ ( .D(n9731), .CLK(clk), .Q(arr[1429]) );
  DFFPOSX1 arr_reg_34__34_ ( .D(n9730), .CLK(clk), .Q(arr[1428]) );
  DFFPOSX1 arr_reg_34__33_ ( .D(n9729), .CLK(clk), .Q(arr[1427]) );
  DFFPOSX1 arr_reg_34__32_ ( .D(n9728), .CLK(clk), .Q(arr[1426]) );
  DFFPOSX1 arr_reg_34__31_ ( .D(n9727), .CLK(clk), .Q(arr[1425]) );
  DFFPOSX1 arr_reg_34__30_ ( .D(n9726), .CLK(clk), .Q(arr[1424]) );
  DFFPOSX1 arr_reg_34__29_ ( .D(n9725), .CLK(clk), .Q(arr[1423]) );
  DFFPOSX1 arr_reg_34__28_ ( .D(n9724), .CLK(clk), .Q(arr[1422]) );
  DFFPOSX1 arr_reg_34__27_ ( .D(n9723), .CLK(clk), .Q(arr[1421]) );
  DFFPOSX1 arr_reg_34__26_ ( .D(n9722), .CLK(clk), .Q(arr[1420]) );
  DFFPOSX1 arr_reg_34__25_ ( .D(n9721), .CLK(clk), .Q(arr[1419]) );
  DFFPOSX1 arr_reg_34__24_ ( .D(n9720), .CLK(clk), .Q(arr[1418]) );
  DFFPOSX1 arr_reg_34__23_ ( .D(n9719), .CLK(clk), .Q(arr[1417]) );
  DFFPOSX1 arr_reg_34__22_ ( .D(n9718), .CLK(clk), .Q(arr[1416]) );
  DFFPOSX1 arr_reg_34__21_ ( .D(n9717), .CLK(clk), .Q(arr[1415]) );
  DFFPOSX1 arr_reg_34__20_ ( .D(n9716), .CLK(clk), .Q(arr[1414]) );
  DFFPOSX1 arr_reg_34__19_ ( .D(n9715), .CLK(clk), .Q(arr[1413]) );
  DFFPOSX1 arr_reg_34__18_ ( .D(n9714), .CLK(clk), .Q(arr[1412]) );
  DFFPOSX1 arr_reg_34__17_ ( .D(n9713), .CLK(clk), .Q(arr[1411]) );
  DFFPOSX1 arr_reg_34__16_ ( .D(n9712), .CLK(clk), .Q(arr[1410]) );
  DFFPOSX1 arr_reg_34__15_ ( .D(n9711), .CLK(clk), .Q(arr[1409]) );
  DFFPOSX1 arr_reg_34__14_ ( .D(n9710), .CLK(clk), .Q(arr[1408]) );
  DFFPOSX1 arr_reg_34__13_ ( .D(n9709), .CLK(clk), .Q(arr[1407]) );
  DFFPOSX1 arr_reg_34__12_ ( .D(n9708), .CLK(clk), .Q(arr[1406]) );
  DFFPOSX1 arr_reg_34__11_ ( .D(n9707), .CLK(clk), .Q(arr[1405]) );
  DFFPOSX1 arr_reg_34__10_ ( .D(n9706), .CLK(clk), .Q(arr[1404]) );
  DFFPOSX1 arr_reg_34__9_ ( .D(n9705), .CLK(clk), .Q(arr[1403]) );
  DFFPOSX1 arr_reg_34__8_ ( .D(n9704), .CLK(clk), .Q(arr[1402]) );
  DFFPOSX1 arr_reg_34__7_ ( .D(n9703), .CLK(clk), .Q(arr[1401]) );
  DFFPOSX1 arr_reg_34__6_ ( .D(n9702), .CLK(clk), .Q(arr[1400]) );
  DFFPOSX1 arr_reg_34__5_ ( .D(n9701), .CLK(clk), .Q(arr[1399]) );
  DFFPOSX1 arr_reg_34__4_ ( .D(n9700), .CLK(clk), .Q(arr[1398]) );
  DFFPOSX1 arr_reg_34__3_ ( .D(n9699), .CLK(clk), .Q(arr[1397]) );
  DFFPOSX1 arr_reg_34__2_ ( .D(n9698), .CLK(clk), .Q(arr[1396]) );
  DFFPOSX1 arr_reg_34__1_ ( .D(n9697), .CLK(clk), .Q(arr[1395]) );
  DFFPOSX1 arr_reg_34__0_ ( .D(n9696), .CLK(clk), .Q(arr[1394]) );
  DFFPOSX1 arr_reg_33__40_ ( .D(n9695), .CLK(clk), .Q(arr[1393]) );
  DFFPOSX1 arr_reg_33__39_ ( .D(n9694), .CLK(clk), .Q(arr[1392]) );
  DFFPOSX1 arr_reg_33__38_ ( .D(n9693), .CLK(clk), .Q(arr[1391]) );
  DFFPOSX1 arr_reg_33__37_ ( .D(n9692), .CLK(clk), .Q(arr[1390]) );
  DFFPOSX1 arr_reg_33__36_ ( .D(n9691), .CLK(clk), .Q(arr[1389]) );
  DFFPOSX1 arr_reg_33__35_ ( .D(n9690), .CLK(clk), .Q(arr[1388]) );
  DFFPOSX1 arr_reg_33__34_ ( .D(n9689), .CLK(clk), .Q(arr[1387]) );
  DFFPOSX1 arr_reg_33__33_ ( .D(n9688), .CLK(clk), .Q(arr[1386]) );
  DFFPOSX1 arr_reg_33__32_ ( .D(n9687), .CLK(clk), .Q(arr[1385]) );
  DFFPOSX1 arr_reg_33__31_ ( .D(n9686), .CLK(clk), .Q(arr[1384]) );
  DFFPOSX1 arr_reg_33__30_ ( .D(n9685), .CLK(clk), .Q(arr[1383]) );
  DFFPOSX1 arr_reg_33__29_ ( .D(n9684), .CLK(clk), .Q(arr[1382]) );
  DFFPOSX1 arr_reg_33__28_ ( .D(n9683), .CLK(clk), .Q(arr[1381]) );
  DFFPOSX1 arr_reg_33__27_ ( .D(n9682), .CLK(clk), .Q(arr[1380]) );
  DFFPOSX1 arr_reg_33__26_ ( .D(n9681), .CLK(clk), .Q(arr[1379]) );
  DFFPOSX1 arr_reg_33__25_ ( .D(n9680), .CLK(clk), .Q(arr[1378]) );
  DFFPOSX1 arr_reg_33__24_ ( .D(n9679), .CLK(clk), .Q(arr[1377]) );
  DFFPOSX1 arr_reg_33__23_ ( .D(n9678), .CLK(clk), .Q(arr[1376]) );
  DFFPOSX1 arr_reg_33__22_ ( .D(n9677), .CLK(clk), .Q(arr[1375]) );
  DFFPOSX1 arr_reg_33__21_ ( .D(n9676), .CLK(clk), .Q(arr[1374]) );
  DFFPOSX1 arr_reg_33__20_ ( .D(n9675), .CLK(clk), .Q(arr[1373]) );
  DFFPOSX1 arr_reg_33__19_ ( .D(n9674), .CLK(clk), .Q(arr[1372]) );
  DFFPOSX1 arr_reg_33__18_ ( .D(n9673), .CLK(clk), .Q(arr[1371]) );
  DFFPOSX1 arr_reg_33__17_ ( .D(n9672), .CLK(clk), .Q(arr[1370]) );
  DFFPOSX1 arr_reg_33__16_ ( .D(n9671), .CLK(clk), .Q(arr[1369]) );
  DFFPOSX1 arr_reg_33__15_ ( .D(n9670), .CLK(clk), .Q(arr[1368]) );
  DFFPOSX1 arr_reg_33__14_ ( .D(n9669), .CLK(clk), .Q(arr[1367]) );
  DFFPOSX1 arr_reg_33__13_ ( .D(n9668), .CLK(clk), .Q(arr[1366]) );
  DFFPOSX1 arr_reg_33__12_ ( .D(n9667), .CLK(clk), .Q(arr[1365]) );
  DFFPOSX1 arr_reg_33__11_ ( .D(n9666), .CLK(clk), .Q(arr[1364]) );
  DFFPOSX1 arr_reg_33__10_ ( .D(n9665), .CLK(clk), .Q(arr[1363]) );
  DFFPOSX1 arr_reg_33__9_ ( .D(n9664), .CLK(clk), .Q(arr[1362]) );
  DFFPOSX1 arr_reg_33__8_ ( .D(n9663), .CLK(clk), .Q(arr[1361]) );
  DFFPOSX1 arr_reg_33__7_ ( .D(n9662), .CLK(clk), .Q(arr[1360]) );
  DFFPOSX1 arr_reg_33__6_ ( .D(n9661), .CLK(clk), .Q(arr[1359]) );
  DFFPOSX1 arr_reg_33__5_ ( .D(n9660), .CLK(clk), .Q(arr[1358]) );
  DFFPOSX1 arr_reg_33__4_ ( .D(n9659), .CLK(clk), .Q(arr[1357]) );
  DFFPOSX1 arr_reg_33__3_ ( .D(n9658), .CLK(clk), .Q(arr[1356]) );
  DFFPOSX1 arr_reg_33__2_ ( .D(n9657), .CLK(clk), .Q(arr[1355]) );
  DFFPOSX1 arr_reg_33__1_ ( .D(n9656), .CLK(clk), .Q(arr[1354]) );
  DFFPOSX1 arr_reg_33__0_ ( .D(n9655), .CLK(clk), .Q(arr[1353]) );
  DFFPOSX1 arr_reg_32__40_ ( .D(n9654), .CLK(clk), .Q(arr[1352]) );
  DFFPOSX1 arr_reg_32__39_ ( .D(n9653), .CLK(clk), .Q(arr[1351]) );
  DFFPOSX1 arr_reg_32__38_ ( .D(n9652), .CLK(clk), .Q(arr[1350]) );
  DFFPOSX1 arr_reg_32__37_ ( .D(n9651), .CLK(clk), .Q(arr[1349]) );
  DFFPOSX1 arr_reg_32__36_ ( .D(n9650), .CLK(clk), .Q(arr[1348]) );
  DFFPOSX1 arr_reg_32__35_ ( .D(n9649), .CLK(clk), .Q(arr[1347]) );
  DFFPOSX1 arr_reg_32__34_ ( .D(n9648), .CLK(clk), .Q(arr[1346]) );
  DFFPOSX1 arr_reg_32__33_ ( .D(n9647), .CLK(clk), .Q(arr[1345]) );
  DFFPOSX1 arr_reg_32__32_ ( .D(n9646), .CLK(clk), .Q(arr[1344]) );
  DFFPOSX1 arr_reg_32__31_ ( .D(n9645), .CLK(clk), .Q(arr[1343]) );
  DFFPOSX1 arr_reg_32__30_ ( .D(n9644), .CLK(clk), .Q(arr[1342]) );
  DFFPOSX1 arr_reg_32__29_ ( .D(n9643), .CLK(clk), .Q(arr[1341]) );
  DFFPOSX1 arr_reg_32__28_ ( .D(n9642), .CLK(clk), .Q(arr[1340]) );
  DFFPOSX1 arr_reg_32__27_ ( .D(n9641), .CLK(clk), .Q(arr[1339]) );
  DFFPOSX1 arr_reg_32__26_ ( .D(n9640), .CLK(clk), .Q(arr[1338]) );
  DFFPOSX1 arr_reg_32__25_ ( .D(n9639), .CLK(clk), .Q(arr[1337]) );
  DFFPOSX1 arr_reg_32__24_ ( .D(n9638), .CLK(clk), .Q(arr[1336]) );
  DFFPOSX1 arr_reg_32__23_ ( .D(n9637), .CLK(clk), .Q(arr[1335]) );
  DFFPOSX1 arr_reg_32__22_ ( .D(n9636), .CLK(clk), .Q(arr[1334]) );
  DFFPOSX1 arr_reg_32__21_ ( .D(n9635), .CLK(clk), .Q(arr[1333]) );
  DFFPOSX1 arr_reg_32__20_ ( .D(n9634), .CLK(clk), .Q(arr[1332]) );
  DFFPOSX1 arr_reg_32__19_ ( .D(n9633), .CLK(clk), .Q(arr[1331]) );
  DFFPOSX1 arr_reg_32__18_ ( .D(n9632), .CLK(clk), .Q(arr[1330]) );
  DFFPOSX1 arr_reg_32__17_ ( .D(n9631), .CLK(clk), .Q(arr[1329]) );
  DFFPOSX1 arr_reg_32__16_ ( .D(n9630), .CLK(clk), .Q(arr[1328]) );
  DFFPOSX1 arr_reg_32__15_ ( .D(n9629), .CLK(clk), .Q(arr[1327]) );
  DFFPOSX1 arr_reg_32__14_ ( .D(n9628), .CLK(clk), .Q(arr[1326]) );
  DFFPOSX1 arr_reg_32__13_ ( .D(n9627), .CLK(clk), .Q(arr[1325]) );
  DFFPOSX1 arr_reg_32__12_ ( .D(n9626), .CLK(clk), .Q(arr[1324]) );
  DFFPOSX1 arr_reg_32__11_ ( .D(n9625), .CLK(clk), .Q(arr[1323]) );
  DFFPOSX1 arr_reg_32__10_ ( .D(n9624), .CLK(clk), .Q(arr[1322]) );
  DFFPOSX1 arr_reg_32__9_ ( .D(n9623), .CLK(clk), .Q(arr[1321]) );
  DFFPOSX1 arr_reg_32__8_ ( .D(n9622), .CLK(clk), .Q(arr[1320]) );
  DFFPOSX1 arr_reg_32__7_ ( .D(n9621), .CLK(clk), .Q(arr[1319]) );
  DFFPOSX1 arr_reg_32__6_ ( .D(n9620), .CLK(clk), .Q(arr[1318]) );
  DFFPOSX1 arr_reg_32__5_ ( .D(n9619), .CLK(clk), .Q(arr[1317]) );
  DFFPOSX1 arr_reg_32__4_ ( .D(n9618), .CLK(clk), .Q(arr[1316]) );
  DFFPOSX1 arr_reg_32__3_ ( .D(n9617), .CLK(clk), .Q(arr[1315]) );
  DFFPOSX1 arr_reg_32__2_ ( .D(n9616), .CLK(clk), .Q(arr[1314]) );
  DFFPOSX1 arr_reg_32__1_ ( .D(n9615), .CLK(clk), .Q(arr[1313]) );
  DFFPOSX1 arr_reg_32__0_ ( .D(n9614), .CLK(clk), .Q(arr[1312]) );
  DFFPOSX1 arr_reg_31__40_ ( .D(n9613), .CLK(clk), .Q(arr[1311]) );
  DFFPOSX1 arr_reg_31__39_ ( .D(n9612), .CLK(clk), .Q(arr[1310]) );
  DFFPOSX1 arr_reg_31__38_ ( .D(n9611), .CLK(clk), .Q(arr[1309]) );
  DFFPOSX1 arr_reg_31__37_ ( .D(n9610), .CLK(clk), .Q(arr[1308]) );
  DFFPOSX1 arr_reg_31__36_ ( .D(n9609), .CLK(clk), .Q(arr[1307]) );
  DFFPOSX1 arr_reg_31__35_ ( .D(n9608), .CLK(clk), .Q(arr[1306]) );
  DFFPOSX1 arr_reg_31__34_ ( .D(n9607), .CLK(clk), .Q(arr[1305]) );
  DFFPOSX1 arr_reg_31__33_ ( .D(n9606), .CLK(clk), .Q(arr[1304]) );
  DFFPOSX1 arr_reg_31__32_ ( .D(n9605), .CLK(clk), .Q(arr[1303]) );
  DFFPOSX1 arr_reg_31__31_ ( .D(n9604), .CLK(clk), .Q(arr[1302]) );
  DFFPOSX1 arr_reg_31__30_ ( .D(n9603), .CLK(clk), .Q(arr[1301]) );
  DFFPOSX1 arr_reg_31__29_ ( .D(n9602), .CLK(clk), .Q(arr[1300]) );
  DFFPOSX1 arr_reg_31__28_ ( .D(n9601), .CLK(clk), .Q(arr[1299]) );
  DFFPOSX1 arr_reg_31__27_ ( .D(n9600), .CLK(clk), .Q(arr[1298]) );
  DFFPOSX1 arr_reg_31__26_ ( .D(n9599), .CLK(clk), .Q(arr[1297]) );
  DFFPOSX1 arr_reg_31__25_ ( .D(n9598), .CLK(clk), .Q(arr[1296]) );
  DFFPOSX1 arr_reg_31__24_ ( .D(n9597), .CLK(clk), .Q(arr[1295]) );
  DFFPOSX1 arr_reg_31__23_ ( .D(n9596), .CLK(clk), .Q(arr[1294]) );
  DFFPOSX1 arr_reg_31__22_ ( .D(n9595), .CLK(clk), .Q(arr[1293]) );
  DFFPOSX1 arr_reg_31__21_ ( .D(n9594), .CLK(clk), .Q(arr[1292]) );
  DFFPOSX1 arr_reg_31__20_ ( .D(n9593), .CLK(clk), .Q(arr[1291]) );
  DFFPOSX1 arr_reg_31__19_ ( .D(n9592), .CLK(clk), .Q(arr[1290]) );
  DFFPOSX1 arr_reg_31__18_ ( .D(n9591), .CLK(clk), .Q(arr[1289]) );
  DFFPOSX1 arr_reg_31__17_ ( .D(n9590), .CLK(clk), .Q(arr[1288]) );
  DFFPOSX1 arr_reg_31__16_ ( .D(n9589), .CLK(clk), .Q(arr[1287]) );
  DFFPOSX1 arr_reg_31__15_ ( .D(n9588), .CLK(clk), .Q(arr[1286]) );
  DFFPOSX1 arr_reg_31__14_ ( .D(n9587), .CLK(clk), .Q(arr[1285]) );
  DFFPOSX1 arr_reg_31__13_ ( .D(n9586), .CLK(clk), .Q(arr[1284]) );
  DFFPOSX1 arr_reg_31__12_ ( .D(n9585), .CLK(clk), .Q(arr[1283]) );
  DFFPOSX1 arr_reg_31__11_ ( .D(n9584), .CLK(clk), .Q(arr[1282]) );
  DFFPOSX1 arr_reg_31__10_ ( .D(n9583), .CLK(clk), .Q(arr[1281]) );
  DFFPOSX1 arr_reg_31__9_ ( .D(n9582), .CLK(clk), .Q(arr[1280]) );
  DFFPOSX1 arr_reg_31__8_ ( .D(n9581), .CLK(clk), .Q(arr[1279]) );
  DFFPOSX1 arr_reg_31__7_ ( .D(n9580), .CLK(clk), .Q(arr[1278]) );
  DFFPOSX1 arr_reg_31__6_ ( .D(n9579), .CLK(clk), .Q(arr[1277]) );
  DFFPOSX1 arr_reg_31__5_ ( .D(n9578), .CLK(clk), .Q(arr[1276]) );
  DFFPOSX1 arr_reg_31__4_ ( .D(n9577), .CLK(clk), .Q(arr[1275]) );
  DFFPOSX1 arr_reg_31__3_ ( .D(n9576), .CLK(clk), .Q(arr[1274]) );
  DFFPOSX1 arr_reg_31__2_ ( .D(n9575), .CLK(clk), .Q(arr[1273]) );
  DFFPOSX1 arr_reg_31__1_ ( .D(n9574), .CLK(clk), .Q(arr[1272]) );
  DFFPOSX1 arr_reg_31__0_ ( .D(n9573), .CLK(clk), .Q(arr[1271]) );
  DFFPOSX1 arr_reg_30__40_ ( .D(n9572), .CLK(clk), .Q(arr[1270]) );
  DFFPOSX1 arr_reg_30__39_ ( .D(n9571), .CLK(clk), .Q(arr[1269]) );
  DFFPOSX1 arr_reg_30__38_ ( .D(n9570), .CLK(clk), .Q(arr[1268]) );
  DFFPOSX1 arr_reg_30__37_ ( .D(n9569), .CLK(clk), .Q(arr[1267]) );
  DFFPOSX1 arr_reg_30__36_ ( .D(n9568), .CLK(clk), .Q(arr[1266]) );
  DFFPOSX1 arr_reg_30__35_ ( .D(n9567), .CLK(clk), .Q(arr[1265]) );
  DFFPOSX1 arr_reg_30__34_ ( .D(n9566), .CLK(clk), .Q(arr[1264]) );
  DFFPOSX1 arr_reg_30__33_ ( .D(n9565), .CLK(clk), .Q(arr[1263]) );
  DFFPOSX1 arr_reg_30__32_ ( .D(n9564), .CLK(clk), .Q(arr[1262]) );
  DFFPOSX1 arr_reg_30__31_ ( .D(n9563), .CLK(clk), .Q(arr[1261]) );
  DFFPOSX1 arr_reg_30__30_ ( .D(n9562), .CLK(clk), .Q(arr[1260]) );
  DFFPOSX1 arr_reg_30__29_ ( .D(n9561), .CLK(clk), .Q(arr[1259]) );
  DFFPOSX1 arr_reg_30__28_ ( .D(n9560), .CLK(clk), .Q(arr[1258]) );
  DFFPOSX1 arr_reg_30__27_ ( .D(n9559), .CLK(clk), .Q(arr[1257]) );
  DFFPOSX1 arr_reg_30__26_ ( .D(n9558), .CLK(clk), .Q(arr[1256]) );
  DFFPOSX1 arr_reg_30__25_ ( .D(n9557), .CLK(clk), .Q(arr[1255]) );
  DFFPOSX1 arr_reg_30__24_ ( .D(n9556), .CLK(clk), .Q(arr[1254]) );
  DFFPOSX1 arr_reg_30__23_ ( .D(n9555), .CLK(clk), .Q(arr[1253]) );
  DFFPOSX1 arr_reg_30__22_ ( .D(n9554), .CLK(clk), .Q(arr[1252]) );
  DFFPOSX1 arr_reg_30__21_ ( .D(n9553), .CLK(clk), .Q(arr[1251]) );
  DFFPOSX1 arr_reg_30__20_ ( .D(n9552), .CLK(clk), .Q(arr[1250]) );
  DFFPOSX1 arr_reg_30__19_ ( .D(n9551), .CLK(clk), .Q(arr[1249]) );
  DFFPOSX1 arr_reg_30__18_ ( .D(n9550), .CLK(clk), .Q(arr[1248]) );
  DFFPOSX1 arr_reg_30__17_ ( .D(n9549), .CLK(clk), .Q(arr[1247]) );
  DFFPOSX1 arr_reg_30__16_ ( .D(n9548), .CLK(clk), .Q(arr[1246]) );
  DFFPOSX1 arr_reg_30__15_ ( .D(n9547), .CLK(clk), .Q(arr[1245]) );
  DFFPOSX1 arr_reg_30__14_ ( .D(n9546), .CLK(clk), .Q(arr[1244]) );
  DFFPOSX1 arr_reg_30__13_ ( .D(n9545), .CLK(clk), .Q(arr[1243]) );
  DFFPOSX1 arr_reg_30__12_ ( .D(n9544), .CLK(clk), .Q(arr[1242]) );
  DFFPOSX1 arr_reg_30__11_ ( .D(n9543), .CLK(clk), .Q(arr[1241]) );
  DFFPOSX1 arr_reg_30__10_ ( .D(n9542), .CLK(clk), .Q(arr[1240]) );
  DFFPOSX1 arr_reg_30__9_ ( .D(n9541), .CLK(clk), .Q(arr[1239]) );
  DFFPOSX1 arr_reg_30__8_ ( .D(n9540), .CLK(clk), .Q(arr[1238]) );
  DFFPOSX1 arr_reg_30__7_ ( .D(n9539), .CLK(clk), .Q(arr[1237]) );
  DFFPOSX1 arr_reg_30__6_ ( .D(n9538), .CLK(clk), .Q(arr[1236]) );
  DFFPOSX1 arr_reg_30__5_ ( .D(n9537), .CLK(clk), .Q(arr[1235]) );
  DFFPOSX1 arr_reg_30__4_ ( .D(n9536), .CLK(clk), .Q(arr[1234]) );
  DFFPOSX1 arr_reg_30__3_ ( .D(n9535), .CLK(clk), .Q(arr[1233]) );
  DFFPOSX1 arr_reg_30__2_ ( .D(n9534), .CLK(clk), .Q(arr[1232]) );
  DFFPOSX1 arr_reg_30__1_ ( .D(n9533), .CLK(clk), .Q(arr[1231]) );
  DFFPOSX1 arr_reg_30__0_ ( .D(n9532), .CLK(clk), .Q(arr[1230]) );
  DFFPOSX1 arr_reg_29__40_ ( .D(n9531), .CLK(clk), .Q(arr[1229]) );
  DFFPOSX1 arr_reg_29__39_ ( .D(n9530), .CLK(clk), .Q(arr[1228]) );
  DFFPOSX1 arr_reg_29__38_ ( .D(n9529), .CLK(clk), .Q(arr[1227]) );
  DFFPOSX1 arr_reg_29__37_ ( .D(n9528), .CLK(clk), .Q(arr[1226]) );
  DFFPOSX1 arr_reg_29__36_ ( .D(n9527), .CLK(clk), .Q(arr[1225]) );
  DFFPOSX1 arr_reg_29__35_ ( .D(n9526), .CLK(clk), .Q(arr[1224]) );
  DFFPOSX1 arr_reg_29__34_ ( .D(n9525), .CLK(clk), .Q(arr[1223]) );
  DFFPOSX1 arr_reg_29__33_ ( .D(n9524), .CLK(clk), .Q(arr[1222]) );
  DFFPOSX1 arr_reg_29__32_ ( .D(n9523), .CLK(clk), .Q(arr[1221]) );
  DFFPOSX1 arr_reg_29__31_ ( .D(n9522), .CLK(clk), .Q(arr[1220]) );
  DFFPOSX1 arr_reg_29__30_ ( .D(n9521), .CLK(clk), .Q(arr[1219]) );
  DFFPOSX1 arr_reg_29__29_ ( .D(n9520), .CLK(clk), .Q(arr[1218]) );
  DFFPOSX1 arr_reg_29__28_ ( .D(n9519), .CLK(clk), .Q(arr[1217]) );
  DFFPOSX1 arr_reg_29__27_ ( .D(n9518), .CLK(clk), .Q(arr[1216]) );
  DFFPOSX1 arr_reg_29__26_ ( .D(n9517), .CLK(clk), .Q(arr[1215]) );
  DFFPOSX1 arr_reg_29__25_ ( .D(n9516), .CLK(clk), .Q(arr[1214]) );
  DFFPOSX1 arr_reg_29__24_ ( .D(n9515), .CLK(clk), .Q(arr[1213]) );
  DFFPOSX1 arr_reg_29__23_ ( .D(n9514), .CLK(clk), .Q(arr[1212]) );
  DFFPOSX1 arr_reg_29__22_ ( .D(n9513), .CLK(clk), .Q(arr[1211]) );
  DFFPOSX1 arr_reg_29__21_ ( .D(n9512), .CLK(clk), .Q(arr[1210]) );
  DFFPOSX1 arr_reg_29__20_ ( .D(n9511), .CLK(clk), .Q(arr[1209]) );
  DFFPOSX1 arr_reg_29__19_ ( .D(n9510), .CLK(clk), .Q(arr[1208]) );
  DFFPOSX1 arr_reg_29__18_ ( .D(n9509), .CLK(clk), .Q(arr[1207]) );
  DFFPOSX1 arr_reg_29__17_ ( .D(n9508), .CLK(clk), .Q(arr[1206]) );
  DFFPOSX1 arr_reg_29__16_ ( .D(n9507), .CLK(clk), .Q(arr[1205]) );
  DFFPOSX1 arr_reg_29__15_ ( .D(n9506), .CLK(clk), .Q(arr[1204]) );
  DFFPOSX1 arr_reg_29__14_ ( .D(n9505), .CLK(clk), .Q(arr[1203]) );
  DFFPOSX1 arr_reg_29__13_ ( .D(n9504), .CLK(clk), .Q(arr[1202]) );
  DFFPOSX1 arr_reg_29__12_ ( .D(n9503), .CLK(clk), .Q(arr[1201]) );
  DFFPOSX1 arr_reg_29__11_ ( .D(n9502), .CLK(clk), .Q(arr[1200]) );
  DFFPOSX1 arr_reg_29__10_ ( .D(n9501), .CLK(clk), .Q(arr[1199]) );
  DFFPOSX1 arr_reg_29__9_ ( .D(n9500), .CLK(clk), .Q(arr[1198]) );
  DFFPOSX1 arr_reg_29__8_ ( .D(n9499), .CLK(clk), .Q(arr[1197]) );
  DFFPOSX1 arr_reg_29__7_ ( .D(n9498), .CLK(clk), .Q(arr[1196]) );
  DFFPOSX1 arr_reg_29__6_ ( .D(n9497), .CLK(clk), .Q(arr[1195]) );
  DFFPOSX1 arr_reg_29__5_ ( .D(n9496), .CLK(clk), .Q(arr[1194]) );
  DFFPOSX1 arr_reg_29__4_ ( .D(n9495), .CLK(clk), .Q(arr[1193]) );
  DFFPOSX1 arr_reg_29__3_ ( .D(n9494), .CLK(clk), .Q(arr[1192]) );
  DFFPOSX1 arr_reg_29__2_ ( .D(n9493), .CLK(clk), .Q(arr[1191]) );
  DFFPOSX1 arr_reg_29__1_ ( .D(n9492), .CLK(clk), .Q(arr[1190]) );
  DFFPOSX1 arr_reg_29__0_ ( .D(n9491), .CLK(clk), .Q(arr[1189]) );
  DFFPOSX1 arr_reg_28__40_ ( .D(n9490), .CLK(clk), .Q(arr[1188]) );
  DFFPOSX1 arr_reg_28__39_ ( .D(n9489), .CLK(clk), .Q(arr[1187]) );
  DFFPOSX1 arr_reg_28__38_ ( .D(n9488), .CLK(clk), .Q(arr[1186]) );
  DFFPOSX1 arr_reg_28__37_ ( .D(n9487), .CLK(clk), .Q(arr[1185]) );
  DFFPOSX1 arr_reg_28__36_ ( .D(n9486), .CLK(clk), .Q(arr[1184]) );
  DFFPOSX1 arr_reg_28__35_ ( .D(n9485), .CLK(clk), .Q(arr[1183]) );
  DFFPOSX1 arr_reg_28__34_ ( .D(n9484), .CLK(clk), .Q(arr[1182]) );
  DFFPOSX1 arr_reg_28__33_ ( .D(n9483), .CLK(clk), .Q(arr[1181]) );
  DFFPOSX1 arr_reg_28__32_ ( .D(n9482), .CLK(clk), .Q(arr[1180]) );
  DFFPOSX1 arr_reg_28__31_ ( .D(n9481), .CLK(clk), .Q(arr[1179]) );
  DFFPOSX1 arr_reg_28__30_ ( .D(n9480), .CLK(clk), .Q(arr[1178]) );
  DFFPOSX1 arr_reg_28__29_ ( .D(n9479), .CLK(clk), .Q(arr[1177]) );
  DFFPOSX1 arr_reg_28__28_ ( .D(n9478), .CLK(clk), .Q(arr[1176]) );
  DFFPOSX1 arr_reg_28__27_ ( .D(n9477), .CLK(clk), .Q(arr[1175]) );
  DFFPOSX1 arr_reg_28__26_ ( .D(n9476), .CLK(clk), .Q(arr[1174]) );
  DFFPOSX1 arr_reg_28__25_ ( .D(n9475), .CLK(clk), .Q(arr[1173]) );
  DFFPOSX1 arr_reg_28__24_ ( .D(n9474), .CLK(clk), .Q(arr[1172]) );
  DFFPOSX1 arr_reg_28__23_ ( .D(n9473), .CLK(clk), .Q(arr[1171]) );
  DFFPOSX1 arr_reg_28__22_ ( .D(n9472), .CLK(clk), .Q(arr[1170]) );
  DFFPOSX1 arr_reg_28__21_ ( .D(n9471), .CLK(clk), .Q(arr[1169]) );
  DFFPOSX1 arr_reg_28__20_ ( .D(n9470), .CLK(clk), .Q(arr[1168]) );
  DFFPOSX1 arr_reg_28__19_ ( .D(n9469), .CLK(clk), .Q(arr[1167]) );
  DFFPOSX1 arr_reg_28__18_ ( .D(n9468), .CLK(clk), .Q(arr[1166]) );
  DFFPOSX1 arr_reg_28__17_ ( .D(n9467), .CLK(clk), .Q(arr[1165]) );
  DFFPOSX1 arr_reg_28__16_ ( .D(n9466), .CLK(clk), .Q(arr[1164]) );
  DFFPOSX1 arr_reg_28__15_ ( .D(n9465), .CLK(clk), .Q(arr[1163]) );
  DFFPOSX1 arr_reg_28__14_ ( .D(n9464), .CLK(clk), .Q(arr[1162]) );
  DFFPOSX1 arr_reg_28__13_ ( .D(n9463), .CLK(clk), .Q(arr[1161]) );
  DFFPOSX1 arr_reg_28__12_ ( .D(n9462), .CLK(clk), .Q(arr[1160]) );
  DFFPOSX1 arr_reg_28__11_ ( .D(n9461), .CLK(clk), .Q(arr[1159]) );
  DFFPOSX1 arr_reg_28__10_ ( .D(n9460), .CLK(clk), .Q(arr[1158]) );
  DFFPOSX1 arr_reg_28__9_ ( .D(n9459), .CLK(clk), .Q(arr[1157]) );
  DFFPOSX1 arr_reg_28__8_ ( .D(n9458), .CLK(clk), .Q(arr[1156]) );
  DFFPOSX1 arr_reg_28__7_ ( .D(n9457), .CLK(clk), .Q(arr[1155]) );
  DFFPOSX1 arr_reg_28__6_ ( .D(n9456), .CLK(clk), .Q(arr[1154]) );
  DFFPOSX1 arr_reg_28__5_ ( .D(n9455), .CLK(clk), .Q(arr[1153]) );
  DFFPOSX1 arr_reg_28__4_ ( .D(n9454), .CLK(clk), .Q(arr[1152]) );
  DFFPOSX1 arr_reg_28__3_ ( .D(n9453), .CLK(clk), .Q(arr[1151]) );
  DFFPOSX1 arr_reg_28__2_ ( .D(n9452), .CLK(clk), .Q(arr[1150]) );
  DFFPOSX1 arr_reg_28__1_ ( .D(n9451), .CLK(clk), .Q(arr[1149]) );
  DFFPOSX1 arr_reg_28__0_ ( .D(n9450), .CLK(clk), .Q(arr[1148]) );
  DFFPOSX1 arr_reg_27__40_ ( .D(n9449), .CLK(clk), .Q(arr[1147]) );
  DFFPOSX1 arr_reg_27__39_ ( .D(n9448), .CLK(clk), .Q(arr[1146]) );
  DFFPOSX1 arr_reg_27__38_ ( .D(n9447), .CLK(clk), .Q(arr[1145]) );
  DFFPOSX1 arr_reg_27__37_ ( .D(n9446), .CLK(clk), .Q(arr[1144]) );
  DFFPOSX1 arr_reg_27__36_ ( .D(n9445), .CLK(clk), .Q(arr[1143]) );
  DFFPOSX1 arr_reg_27__35_ ( .D(n9444), .CLK(clk), .Q(arr[1142]) );
  DFFPOSX1 arr_reg_27__34_ ( .D(n9443), .CLK(clk), .Q(arr[1141]) );
  DFFPOSX1 arr_reg_27__33_ ( .D(n9442), .CLK(clk), .Q(arr[1140]) );
  DFFPOSX1 arr_reg_27__32_ ( .D(n9441), .CLK(clk), .Q(arr[1139]) );
  DFFPOSX1 arr_reg_27__31_ ( .D(n9440), .CLK(clk), .Q(arr[1138]) );
  DFFPOSX1 arr_reg_27__30_ ( .D(n9439), .CLK(clk), .Q(arr[1137]) );
  DFFPOSX1 arr_reg_27__29_ ( .D(n9438), .CLK(clk), .Q(arr[1136]) );
  DFFPOSX1 arr_reg_27__28_ ( .D(n9437), .CLK(clk), .Q(arr[1135]) );
  DFFPOSX1 arr_reg_27__27_ ( .D(n9436), .CLK(clk), .Q(arr[1134]) );
  DFFPOSX1 arr_reg_27__26_ ( .D(n9435), .CLK(clk), .Q(arr[1133]) );
  DFFPOSX1 arr_reg_27__25_ ( .D(n9434), .CLK(clk), .Q(arr[1132]) );
  DFFPOSX1 arr_reg_27__24_ ( .D(n9433), .CLK(clk), .Q(arr[1131]) );
  DFFPOSX1 arr_reg_27__23_ ( .D(n9432), .CLK(clk), .Q(arr[1130]) );
  DFFPOSX1 arr_reg_27__22_ ( .D(n9431), .CLK(clk), .Q(arr[1129]) );
  DFFPOSX1 arr_reg_27__21_ ( .D(n9430), .CLK(clk), .Q(arr[1128]) );
  DFFPOSX1 arr_reg_27__20_ ( .D(n9429), .CLK(clk), .Q(arr[1127]) );
  DFFPOSX1 arr_reg_27__19_ ( .D(n9428), .CLK(clk), .Q(arr[1126]) );
  DFFPOSX1 arr_reg_27__18_ ( .D(n9427), .CLK(clk), .Q(arr[1125]) );
  DFFPOSX1 arr_reg_27__17_ ( .D(n9426), .CLK(clk), .Q(arr[1124]) );
  DFFPOSX1 arr_reg_27__16_ ( .D(n9425), .CLK(clk), .Q(arr[1123]) );
  DFFPOSX1 arr_reg_27__15_ ( .D(n9424), .CLK(clk), .Q(arr[1122]) );
  DFFPOSX1 arr_reg_27__14_ ( .D(n9423), .CLK(clk), .Q(arr[1121]) );
  DFFPOSX1 arr_reg_27__13_ ( .D(n9422), .CLK(clk), .Q(arr[1120]) );
  DFFPOSX1 arr_reg_27__12_ ( .D(n9421), .CLK(clk), .Q(arr[1119]) );
  DFFPOSX1 arr_reg_27__11_ ( .D(n9420), .CLK(clk), .Q(arr[1118]) );
  DFFPOSX1 arr_reg_27__10_ ( .D(n9419), .CLK(clk), .Q(arr[1117]) );
  DFFPOSX1 arr_reg_27__9_ ( .D(n9418), .CLK(clk), .Q(arr[1116]) );
  DFFPOSX1 arr_reg_27__8_ ( .D(n9417), .CLK(clk), .Q(arr[1115]) );
  DFFPOSX1 arr_reg_27__7_ ( .D(n9416), .CLK(clk), .Q(arr[1114]) );
  DFFPOSX1 arr_reg_27__6_ ( .D(n9415), .CLK(clk), .Q(arr[1113]) );
  DFFPOSX1 arr_reg_27__5_ ( .D(n9414), .CLK(clk), .Q(arr[1112]) );
  DFFPOSX1 arr_reg_27__4_ ( .D(n9413), .CLK(clk), .Q(arr[1111]) );
  DFFPOSX1 arr_reg_27__3_ ( .D(n9412), .CLK(clk), .Q(arr[1110]) );
  DFFPOSX1 arr_reg_27__2_ ( .D(n9411), .CLK(clk), .Q(arr[1109]) );
  DFFPOSX1 arr_reg_27__1_ ( .D(n9410), .CLK(clk), .Q(arr[1108]) );
  DFFPOSX1 arr_reg_27__0_ ( .D(n9409), .CLK(clk), .Q(arr[1107]) );
  DFFPOSX1 arr_reg_26__40_ ( .D(n9408), .CLK(clk), .Q(arr[1106]) );
  DFFPOSX1 arr_reg_26__39_ ( .D(n9407), .CLK(clk), .Q(arr[1105]) );
  DFFPOSX1 arr_reg_26__38_ ( .D(n9406), .CLK(clk), .Q(arr[1104]) );
  DFFPOSX1 arr_reg_26__37_ ( .D(n9405), .CLK(clk), .Q(arr[1103]) );
  DFFPOSX1 arr_reg_26__36_ ( .D(n9404), .CLK(clk), .Q(arr[1102]) );
  DFFPOSX1 arr_reg_26__35_ ( .D(n9403), .CLK(clk), .Q(arr[1101]) );
  DFFPOSX1 arr_reg_26__34_ ( .D(n9402), .CLK(clk), .Q(arr[1100]) );
  DFFPOSX1 arr_reg_26__33_ ( .D(n9401), .CLK(clk), .Q(arr[1099]) );
  DFFPOSX1 arr_reg_26__32_ ( .D(n9400), .CLK(clk), .Q(arr[1098]) );
  DFFPOSX1 arr_reg_26__31_ ( .D(n9399), .CLK(clk), .Q(arr[1097]) );
  DFFPOSX1 arr_reg_26__30_ ( .D(n9398), .CLK(clk), .Q(arr[1096]) );
  DFFPOSX1 arr_reg_26__29_ ( .D(n9397), .CLK(clk), .Q(arr[1095]) );
  DFFPOSX1 arr_reg_26__28_ ( .D(n9396), .CLK(clk), .Q(arr[1094]) );
  DFFPOSX1 arr_reg_26__27_ ( .D(n9395), .CLK(clk), .Q(arr[1093]) );
  DFFPOSX1 arr_reg_26__26_ ( .D(n9394), .CLK(clk), .Q(arr[1092]) );
  DFFPOSX1 arr_reg_26__25_ ( .D(n9393), .CLK(clk), .Q(arr[1091]) );
  DFFPOSX1 arr_reg_26__24_ ( .D(n9392), .CLK(clk), .Q(arr[1090]) );
  DFFPOSX1 arr_reg_26__23_ ( .D(n9391), .CLK(clk), .Q(arr[1089]) );
  DFFPOSX1 arr_reg_26__22_ ( .D(n9390), .CLK(clk), .Q(arr[1088]) );
  DFFPOSX1 arr_reg_26__21_ ( .D(n9389), .CLK(clk), .Q(arr[1087]) );
  DFFPOSX1 arr_reg_26__20_ ( .D(n9388), .CLK(clk), .Q(arr[1086]) );
  DFFPOSX1 arr_reg_26__19_ ( .D(n9387), .CLK(clk), .Q(arr[1085]) );
  DFFPOSX1 arr_reg_26__18_ ( .D(n9386), .CLK(clk), .Q(arr[1084]) );
  DFFPOSX1 arr_reg_26__17_ ( .D(n9385), .CLK(clk), .Q(arr[1083]) );
  DFFPOSX1 arr_reg_26__16_ ( .D(n9384), .CLK(clk), .Q(arr[1082]) );
  DFFPOSX1 arr_reg_26__15_ ( .D(n9383), .CLK(clk), .Q(arr[1081]) );
  DFFPOSX1 arr_reg_26__14_ ( .D(n9382), .CLK(clk), .Q(arr[1080]) );
  DFFPOSX1 arr_reg_26__13_ ( .D(n9381), .CLK(clk), .Q(arr[1079]) );
  DFFPOSX1 arr_reg_26__12_ ( .D(n9380), .CLK(clk), .Q(arr[1078]) );
  DFFPOSX1 arr_reg_26__11_ ( .D(n9379), .CLK(clk), .Q(arr[1077]) );
  DFFPOSX1 arr_reg_26__10_ ( .D(n9378), .CLK(clk), .Q(arr[1076]) );
  DFFPOSX1 arr_reg_26__9_ ( .D(n9377), .CLK(clk), .Q(arr[1075]) );
  DFFPOSX1 arr_reg_26__8_ ( .D(n9376), .CLK(clk), .Q(arr[1074]) );
  DFFPOSX1 arr_reg_26__7_ ( .D(n9375), .CLK(clk), .Q(arr[1073]) );
  DFFPOSX1 arr_reg_26__6_ ( .D(n9374), .CLK(clk), .Q(arr[1072]) );
  DFFPOSX1 arr_reg_26__5_ ( .D(n9373), .CLK(clk), .Q(arr[1071]) );
  DFFPOSX1 arr_reg_26__4_ ( .D(n9372), .CLK(clk), .Q(arr[1070]) );
  DFFPOSX1 arr_reg_26__3_ ( .D(n9371), .CLK(clk), .Q(arr[1069]) );
  DFFPOSX1 arr_reg_26__2_ ( .D(n9370), .CLK(clk), .Q(arr[1068]) );
  DFFPOSX1 arr_reg_26__1_ ( .D(n9369), .CLK(clk), .Q(arr[1067]) );
  DFFPOSX1 arr_reg_26__0_ ( .D(n9368), .CLK(clk), .Q(arr[1066]) );
  DFFPOSX1 arr_reg_25__40_ ( .D(n9367), .CLK(clk), .Q(arr[1065]) );
  DFFPOSX1 arr_reg_25__39_ ( .D(n9366), .CLK(clk), .Q(arr[1064]) );
  DFFPOSX1 arr_reg_25__38_ ( .D(n9365), .CLK(clk), .Q(arr[1063]) );
  DFFPOSX1 arr_reg_25__37_ ( .D(n9364), .CLK(clk), .Q(arr[1062]) );
  DFFPOSX1 arr_reg_25__36_ ( .D(n9363), .CLK(clk), .Q(arr[1061]) );
  DFFPOSX1 arr_reg_25__35_ ( .D(n9362), .CLK(clk), .Q(arr[1060]) );
  DFFPOSX1 arr_reg_25__34_ ( .D(n9361), .CLK(clk), .Q(arr[1059]) );
  DFFPOSX1 arr_reg_25__33_ ( .D(n9360), .CLK(clk), .Q(arr[1058]) );
  DFFPOSX1 arr_reg_25__32_ ( .D(n9359), .CLK(clk), .Q(arr[1057]) );
  DFFPOSX1 arr_reg_25__31_ ( .D(n9358), .CLK(clk), .Q(arr[1056]) );
  DFFPOSX1 arr_reg_25__30_ ( .D(n9357), .CLK(clk), .Q(arr[1055]) );
  DFFPOSX1 arr_reg_25__29_ ( .D(n9356), .CLK(clk), .Q(arr[1054]) );
  DFFPOSX1 arr_reg_25__28_ ( .D(n9355), .CLK(clk), .Q(arr[1053]) );
  DFFPOSX1 arr_reg_25__27_ ( .D(n9354), .CLK(clk), .Q(arr[1052]) );
  DFFPOSX1 arr_reg_25__26_ ( .D(n9353), .CLK(clk), .Q(arr[1051]) );
  DFFPOSX1 arr_reg_25__25_ ( .D(n9352), .CLK(clk), .Q(arr[1050]) );
  DFFPOSX1 arr_reg_25__24_ ( .D(n9351), .CLK(clk), .Q(arr[1049]) );
  DFFPOSX1 arr_reg_25__23_ ( .D(n9350), .CLK(clk), .Q(arr[1048]) );
  DFFPOSX1 arr_reg_25__22_ ( .D(n9349), .CLK(clk), .Q(arr[1047]) );
  DFFPOSX1 arr_reg_25__21_ ( .D(n9348), .CLK(clk), .Q(arr[1046]) );
  DFFPOSX1 arr_reg_25__20_ ( .D(n9347), .CLK(clk), .Q(arr[1045]) );
  DFFPOSX1 arr_reg_25__19_ ( .D(n9346), .CLK(clk), .Q(arr[1044]) );
  DFFPOSX1 arr_reg_25__18_ ( .D(n9345), .CLK(clk), .Q(arr[1043]) );
  DFFPOSX1 arr_reg_25__17_ ( .D(n9344), .CLK(clk), .Q(arr[1042]) );
  DFFPOSX1 arr_reg_25__16_ ( .D(n9343), .CLK(clk), .Q(arr[1041]) );
  DFFPOSX1 arr_reg_25__15_ ( .D(n9342), .CLK(clk), .Q(arr[1040]) );
  DFFPOSX1 arr_reg_25__14_ ( .D(n9341), .CLK(clk), .Q(arr[1039]) );
  DFFPOSX1 arr_reg_25__13_ ( .D(n9340), .CLK(clk), .Q(arr[1038]) );
  DFFPOSX1 arr_reg_25__12_ ( .D(n9339), .CLK(clk), .Q(arr[1037]) );
  DFFPOSX1 arr_reg_25__11_ ( .D(n9338), .CLK(clk), .Q(arr[1036]) );
  DFFPOSX1 arr_reg_25__10_ ( .D(n9337), .CLK(clk), .Q(arr[1035]) );
  DFFPOSX1 arr_reg_25__9_ ( .D(n9336), .CLK(clk), .Q(arr[1034]) );
  DFFPOSX1 arr_reg_25__8_ ( .D(n9335), .CLK(clk), .Q(arr[1033]) );
  DFFPOSX1 arr_reg_25__7_ ( .D(n9334), .CLK(clk), .Q(arr[1032]) );
  DFFPOSX1 arr_reg_25__6_ ( .D(n9333), .CLK(clk), .Q(arr[1031]) );
  DFFPOSX1 arr_reg_25__5_ ( .D(n9332), .CLK(clk), .Q(arr[1030]) );
  DFFPOSX1 arr_reg_25__4_ ( .D(n9331), .CLK(clk), .Q(arr[1029]) );
  DFFPOSX1 arr_reg_25__3_ ( .D(n9330), .CLK(clk), .Q(arr[1028]) );
  DFFPOSX1 arr_reg_25__2_ ( .D(n9329), .CLK(clk), .Q(arr[1027]) );
  DFFPOSX1 arr_reg_25__1_ ( .D(n9328), .CLK(clk), .Q(arr[1026]) );
  DFFPOSX1 arr_reg_25__0_ ( .D(n9327), .CLK(clk), .Q(arr[1025]) );
  DFFPOSX1 arr_reg_24__40_ ( .D(n9326), .CLK(clk), .Q(arr[1024]) );
  DFFPOSX1 arr_reg_24__39_ ( .D(n9325), .CLK(clk), .Q(arr[1023]) );
  DFFPOSX1 arr_reg_24__38_ ( .D(n9324), .CLK(clk), .Q(arr[1022]) );
  DFFPOSX1 arr_reg_24__37_ ( .D(n9323), .CLK(clk), .Q(arr[1021]) );
  DFFPOSX1 arr_reg_24__36_ ( .D(n9322), .CLK(clk), .Q(arr[1020]) );
  DFFPOSX1 arr_reg_24__35_ ( .D(n9321), .CLK(clk), .Q(arr[1019]) );
  DFFPOSX1 arr_reg_24__34_ ( .D(n9320), .CLK(clk), .Q(arr[1018]) );
  DFFPOSX1 arr_reg_24__33_ ( .D(n9319), .CLK(clk), .Q(arr[1017]) );
  DFFPOSX1 arr_reg_24__32_ ( .D(n9318), .CLK(clk), .Q(arr[1016]) );
  DFFPOSX1 arr_reg_24__31_ ( .D(n9317), .CLK(clk), .Q(arr[1015]) );
  DFFPOSX1 arr_reg_24__30_ ( .D(n9316), .CLK(clk), .Q(arr[1014]) );
  DFFPOSX1 arr_reg_24__29_ ( .D(n9315), .CLK(clk), .Q(arr[1013]) );
  DFFPOSX1 arr_reg_24__28_ ( .D(n9314), .CLK(clk), .Q(arr[1012]) );
  DFFPOSX1 arr_reg_24__27_ ( .D(n9313), .CLK(clk), .Q(arr[1011]) );
  DFFPOSX1 arr_reg_24__26_ ( .D(n9312), .CLK(clk), .Q(arr[1010]) );
  DFFPOSX1 arr_reg_24__25_ ( .D(n9311), .CLK(clk), .Q(arr[1009]) );
  DFFPOSX1 arr_reg_24__24_ ( .D(n9310), .CLK(clk), .Q(arr[1008]) );
  DFFPOSX1 arr_reg_24__23_ ( .D(n9309), .CLK(clk), .Q(arr[1007]) );
  DFFPOSX1 arr_reg_24__22_ ( .D(n9308), .CLK(clk), .Q(arr[1006]) );
  DFFPOSX1 arr_reg_24__21_ ( .D(n9307), .CLK(clk), .Q(arr[1005]) );
  DFFPOSX1 arr_reg_24__20_ ( .D(n9306), .CLK(clk), .Q(arr[1004]) );
  DFFPOSX1 arr_reg_24__19_ ( .D(n9305), .CLK(clk), .Q(arr[1003]) );
  DFFPOSX1 arr_reg_24__18_ ( .D(n9304), .CLK(clk), .Q(arr[1002]) );
  DFFPOSX1 arr_reg_24__17_ ( .D(n9303), .CLK(clk), .Q(arr[1001]) );
  DFFPOSX1 arr_reg_24__16_ ( .D(n9302), .CLK(clk), .Q(arr[1000]) );
  DFFPOSX1 arr_reg_24__15_ ( .D(n9301), .CLK(clk), .Q(arr[999]) );
  DFFPOSX1 arr_reg_24__14_ ( .D(n9300), .CLK(clk), .Q(arr[998]) );
  DFFPOSX1 arr_reg_24__13_ ( .D(n9299), .CLK(clk), .Q(arr[997]) );
  DFFPOSX1 arr_reg_24__12_ ( .D(n9298), .CLK(clk), .Q(arr[996]) );
  DFFPOSX1 arr_reg_24__11_ ( .D(n9297), .CLK(clk), .Q(arr[995]) );
  DFFPOSX1 arr_reg_24__10_ ( .D(n9296), .CLK(clk), .Q(arr[994]) );
  DFFPOSX1 arr_reg_24__9_ ( .D(n9295), .CLK(clk), .Q(arr[993]) );
  DFFPOSX1 arr_reg_24__8_ ( .D(n9294), .CLK(clk), .Q(arr[992]) );
  DFFPOSX1 arr_reg_24__7_ ( .D(n9293), .CLK(clk), .Q(arr[991]) );
  DFFPOSX1 arr_reg_24__6_ ( .D(n9292), .CLK(clk), .Q(arr[990]) );
  DFFPOSX1 arr_reg_24__5_ ( .D(n9291), .CLK(clk), .Q(arr[989]) );
  DFFPOSX1 arr_reg_24__4_ ( .D(n9290), .CLK(clk), .Q(arr[988]) );
  DFFPOSX1 arr_reg_24__3_ ( .D(n9289), .CLK(clk), .Q(arr[987]) );
  DFFPOSX1 arr_reg_24__2_ ( .D(n9288), .CLK(clk), .Q(arr[986]) );
  DFFPOSX1 arr_reg_24__1_ ( .D(n9287), .CLK(clk), .Q(arr[985]) );
  DFFPOSX1 arr_reg_24__0_ ( .D(n9286), .CLK(clk), .Q(arr[984]) );
  DFFPOSX1 arr_reg_23__40_ ( .D(n9285), .CLK(clk), .Q(arr[983]) );
  DFFPOSX1 arr_reg_23__39_ ( .D(n9284), .CLK(clk), .Q(arr[982]) );
  DFFPOSX1 arr_reg_23__38_ ( .D(n9283), .CLK(clk), .Q(arr[981]) );
  DFFPOSX1 arr_reg_23__37_ ( .D(n9282), .CLK(clk), .Q(arr[980]) );
  DFFPOSX1 arr_reg_23__36_ ( .D(n9281), .CLK(clk), .Q(arr[979]) );
  DFFPOSX1 arr_reg_23__35_ ( .D(n9280), .CLK(clk), .Q(arr[978]) );
  DFFPOSX1 arr_reg_23__34_ ( .D(n9279), .CLK(clk), .Q(arr[977]) );
  DFFPOSX1 arr_reg_23__33_ ( .D(n9278), .CLK(clk), .Q(arr[976]) );
  DFFPOSX1 arr_reg_23__32_ ( .D(n9277), .CLK(clk), .Q(arr[975]) );
  DFFPOSX1 arr_reg_23__31_ ( .D(n9276), .CLK(clk), .Q(arr[974]) );
  DFFPOSX1 arr_reg_23__30_ ( .D(n9275), .CLK(clk), .Q(arr[973]) );
  DFFPOSX1 arr_reg_23__29_ ( .D(n9274), .CLK(clk), .Q(arr[972]) );
  DFFPOSX1 arr_reg_23__28_ ( .D(n9273), .CLK(clk), .Q(arr[971]) );
  DFFPOSX1 arr_reg_23__27_ ( .D(n9272), .CLK(clk), .Q(arr[970]) );
  DFFPOSX1 arr_reg_23__26_ ( .D(n9271), .CLK(clk), .Q(arr[969]) );
  DFFPOSX1 arr_reg_23__25_ ( .D(n9270), .CLK(clk), .Q(arr[968]) );
  DFFPOSX1 arr_reg_23__24_ ( .D(n9269), .CLK(clk), .Q(arr[967]) );
  DFFPOSX1 arr_reg_23__23_ ( .D(n9268), .CLK(clk), .Q(arr[966]) );
  DFFPOSX1 arr_reg_23__22_ ( .D(n9267), .CLK(clk), .Q(arr[965]) );
  DFFPOSX1 arr_reg_23__21_ ( .D(n9266), .CLK(clk), .Q(arr[964]) );
  DFFPOSX1 arr_reg_23__20_ ( .D(n9265), .CLK(clk), .Q(arr[963]) );
  DFFPOSX1 arr_reg_23__19_ ( .D(n9264), .CLK(clk), .Q(arr[962]) );
  DFFPOSX1 arr_reg_23__18_ ( .D(n9263), .CLK(clk), .Q(arr[961]) );
  DFFPOSX1 arr_reg_23__17_ ( .D(n9262), .CLK(clk), .Q(arr[960]) );
  DFFPOSX1 arr_reg_23__16_ ( .D(n9261), .CLK(clk), .Q(arr[959]) );
  DFFPOSX1 arr_reg_23__15_ ( .D(n9260), .CLK(clk), .Q(arr[958]) );
  DFFPOSX1 arr_reg_23__14_ ( .D(n9259), .CLK(clk), .Q(arr[957]) );
  DFFPOSX1 arr_reg_23__13_ ( .D(n9258), .CLK(clk), .Q(arr[956]) );
  DFFPOSX1 arr_reg_23__12_ ( .D(n9257), .CLK(clk), .Q(arr[955]) );
  DFFPOSX1 arr_reg_23__11_ ( .D(n9256), .CLK(clk), .Q(arr[954]) );
  DFFPOSX1 arr_reg_23__10_ ( .D(n9255), .CLK(clk), .Q(arr[953]) );
  DFFPOSX1 arr_reg_23__9_ ( .D(n9254), .CLK(clk), .Q(arr[952]) );
  DFFPOSX1 arr_reg_23__8_ ( .D(n9253), .CLK(clk), .Q(arr[951]) );
  DFFPOSX1 arr_reg_23__7_ ( .D(n9252), .CLK(clk), .Q(arr[950]) );
  DFFPOSX1 arr_reg_23__6_ ( .D(n9251), .CLK(clk), .Q(arr[949]) );
  DFFPOSX1 arr_reg_23__5_ ( .D(n9250), .CLK(clk), .Q(arr[948]) );
  DFFPOSX1 arr_reg_23__4_ ( .D(n9249), .CLK(clk), .Q(arr[947]) );
  DFFPOSX1 arr_reg_23__3_ ( .D(n9248), .CLK(clk), .Q(arr[946]) );
  DFFPOSX1 arr_reg_23__2_ ( .D(n9247), .CLK(clk), .Q(arr[945]) );
  DFFPOSX1 arr_reg_23__1_ ( .D(n9246), .CLK(clk), .Q(arr[944]) );
  DFFPOSX1 arr_reg_23__0_ ( .D(n9245), .CLK(clk), .Q(arr[943]) );
  DFFPOSX1 arr_reg_22__40_ ( .D(n9244), .CLK(clk), .Q(arr[942]) );
  DFFPOSX1 arr_reg_22__39_ ( .D(n9243), .CLK(clk), .Q(arr[941]) );
  DFFPOSX1 arr_reg_22__38_ ( .D(n9242), .CLK(clk), .Q(arr[940]) );
  DFFPOSX1 arr_reg_22__37_ ( .D(n9241), .CLK(clk), .Q(arr[939]) );
  DFFPOSX1 arr_reg_22__36_ ( .D(n9240), .CLK(clk), .Q(arr[938]) );
  DFFPOSX1 arr_reg_22__35_ ( .D(n9239), .CLK(clk), .Q(arr[937]) );
  DFFPOSX1 arr_reg_22__34_ ( .D(n9238), .CLK(clk), .Q(arr[936]) );
  DFFPOSX1 arr_reg_22__33_ ( .D(n9237), .CLK(clk), .Q(arr[935]) );
  DFFPOSX1 arr_reg_22__32_ ( .D(n9236), .CLK(clk), .Q(arr[934]) );
  DFFPOSX1 arr_reg_22__31_ ( .D(n9235), .CLK(clk), .Q(arr[933]) );
  DFFPOSX1 arr_reg_22__30_ ( .D(n9234), .CLK(clk), .Q(arr[932]) );
  DFFPOSX1 arr_reg_22__29_ ( .D(n9233), .CLK(clk), .Q(arr[931]) );
  DFFPOSX1 arr_reg_22__28_ ( .D(n9232), .CLK(clk), .Q(arr[930]) );
  DFFPOSX1 arr_reg_22__27_ ( .D(n9231), .CLK(clk), .Q(arr[929]) );
  DFFPOSX1 arr_reg_22__26_ ( .D(n9230), .CLK(clk), .Q(arr[928]) );
  DFFPOSX1 arr_reg_22__25_ ( .D(n9229), .CLK(clk), .Q(arr[927]) );
  DFFPOSX1 arr_reg_22__24_ ( .D(n9228), .CLK(clk), .Q(arr[926]) );
  DFFPOSX1 arr_reg_22__23_ ( .D(n9227), .CLK(clk), .Q(arr[925]) );
  DFFPOSX1 arr_reg_22__22_ ( .D(n9226), .CLK(clk), .Q(arr[924]) );
  DFFPOSX1 arr_reg_22__21_ ( .D(n9225), .CLK(clk), .Q(arr[923]) );
  DFFPOSX1 arr_reg_22__20_ ( .D(n9224), .CLK(clk), .Q(arr[922]) );
  DFFPOSX1 arr_reg_22__19_ ( .D(n9223), .CLK(clk), .Q(arr[921]) );
  DFFPOSX1 arr_reg_22__18_ ( .D(n9222), .CLK(clk), .Q(arr[920]) );
  DFFPOSX1 arr_reg_22__17_ ( .D(n9221), .CLK(clk), .Q(arr[919]) );
  DFFPOSX1 arr_reg_22__16_ ( .D(n9220), .CLK(clk), .Q(arr[918]) );
  DFFPOSX1 arr_reg_22__15_ ( .D(n9219), .CLK(clk), .Q(arr[917]) );
  DFFPOSX1 arr_reg_22__14_ ( .D(n9218), .CLK(clk), .Q(arr[916]) );
  DFFPOSX1 arr_reg_22__13_ ( .D(n9217), .CLK(clk), .Q(arr[915]) );
  DFFPOSX1 arr_reg_22__12_ ( .D(n9216), .CLK(clk), .Q(arr[914]) );
  DFFPOSX1 arr_reg_22__11_ ( .D(n9215), .CLK(clk), .Q(arr[913]) );
  DFFPOSX1 arr_reg_22__10_ ( .D(n9214), .CLK(clk), .Q(arr[912]) );
  DFFPOSX1 arr_reg_22__9_ ( .D(n9213), .CLK(clk), .Q(arr[911]) );
  DFFPOSX1 arr_reg_22__8_ ( .D(n9212), .CLK(clk), .Q(arr[910]) );
  DFFPOSX1 arr_reg_22__7_ ( .D(n9211), .CLK(clk), .Q(arr[909]) );
  DFFPOSX1 arr_reg_22__6_ ( .D(n9210), .CLK(clk), .Q(arr[908]) );
  DFFPOSX1 arr_reg_22__5_ ( .D(n9209), .CLK(clk), .Q(arr[907]) );
  DFFPOSX1 arr_reg_22__4_ ( .D(n9208), .CLK(clk), .Q(arr[906]) );
  DFFPOSX1 arr_reg_22__3_ ( .D(n9207), .CLK(clk), .Q(arr[905]) );
  DFFPOSX1 arr_reg_22__2_ ( .D(n9206), .CLK(clk), .Q(arr[904]) );
  DFFPOSX1 arr_reg_22__1_ ( .D(n9205), .CLK(clk), .Q(arr[903]) );
  DFFPOSX1 arr_reg_22__0_ ( .D(n9204), .CLK(clk), .Q(arr[902]) );
  DFFPOSX1 arr_reg_21__40_ ( .D(n9203), .CLK(clk), .Q(arr[901]) );
  DFFPOSX1 arr_reg_21__39_ ( .D(n9202), .CLK(clk), .Q(arr[900]) );
  DFFPOSX1 arr_reg_21__38_ ( .D(n9201), .CLK(clk), .Q(arr[899]) );
  DFFPOSX1 arr_reg_21__37_ ( .D(n9200), .CLK(clk), .Q(arr[898]) );
  DFFPOSX1 arr_reg_21__36_ ( .D(n9199), .CLK(clk), .Q(arr[897]) );
  DFFPOSX1 arr_reg_21__35_ ( .D(n9198), .CLK(clk), .Q(arr[896]) );
  DFFPOSX1 arr_reg_21__34_ ( .D(n9197), .CLK(clk), .Q(arr[895]) );
  DFFPOSX1 arr_reg_21__33_ ( .D(n9196), .CLK(clk), .Q(arr[894]) );
  DFFPOSX1 arr_reg_21__32_ ( .D(n9195), .CLK(clk), .Q(arr[893]) );
  DFFPOSX1 arr_reg_21__31_ ( .D(n9194), .CLK(clk), .Q(arr[892]) );
  DFFPOSX1 arr_reg_21__30_ ( .D(n9193), .CLK(clk), .Q(arr[891]) );
  DFFPOSX1 arr_reg_21__29_ ( .D(n9192), .CLK(clk), .Q(arr[890]) );
  DFFPOSX1 arr_reg_21__28_ ( .D(n9191), .CLK(clk), .Q(arr[889]) );
  DFFPOSX1 arr_reg_21__27_ ( .D(n9190), .CLK(clk), .Q(arr[888]) );
  DFFPOSX1 arr_reg_21__26_ ( .D(n9189), .CLK(clk), .Q(arr[887]) );
  DFFPOSX1 arr_reg_21__25_ ( .D(n9188), .CLK(clk), .Q(arr[886]) );
  DFFPOSX1 arr_reg_21__24_ ( .D(n9187), .CLK(clk), .Q(arr[885]) );
  DFFPOSX1 arr_reg_21__23_ ( .D(n9186), .CLK(clk), .Q(arr[884]) );
  DFFPOSX1 arr_reg_21__22_ ( .D(n9185), .CLK(clk), .Q(arr[883]) );
  DFFPOSX1 arr_reg_21__21_ ( .D(n9184), .CLK(clk), .Q(arr[882]) );
  DFFPOSX1 arr_reg_21__20_ ( .D(n9183), .CLK(clk), .Q(arr[881]) );
  DFFPOSX1 arr_reg_21__19_ ( .D(n9182), .CLK(clk), .Q(arr[880]) );
  DFFPOSX1 arr_reg_21__18_ ( .D(n9181), .CLK(clk), .Q(arr[879]) );
  DFFPOSX1 arr_reg_21__17_ ( .D(n9180), .CLK(clk), .Q(arr[878]) );
  DFFPOSX1 arr_reg_21__16_ ( .D(n9179), .CLK(clk), .Q(arr[877]) );
  DFFPOSX1 arr_reg_21__15_ ( .D(n9178), .CLK(clk), .Q(arr[876]) );
  DFFPOSX1 arr_reg_21__14_ ( .D(n9177), .CLK(clk), .Q(arr[875]) );
  DFFPOSX1 arr_reg_21__13_ ( .D(n9176), .CLK(clk), .Q(arr[874]) );
  DFFPOSX1 arr_reg_21__12_ ( .D(n9175), .CLK(clk), .Q(arr[873]) );
  DFFPOSX1 arr_reg_21__11_ ( .D(n9174), .CLK(clk), .Q(arr[872]) );
  DFFPOSX1 arr_reg_21__10_ ( .D(n9173), .CLK(clk), .Q(arr[871]) );
  DFFPOSX1 arr_reg_21__9_ ( .D(n9172), .CLK(clk), .Q(arr[870]) );
  DFFPOSX1 arr_reg_21__8_ ( .D(n9171), .CLK(clk), .Q(arr[869]) );
  DFFPOSX1 arr_reg_21__7_ ( .D(n9170), .CLK(clk), .Q(arr[868]) );
  DFFPOSX1 arr_reg_21__6_ ( .D(n9169), .CLK(clk), .Q(arr[867]) );
  DFFPOSX1 arr_reg_21__5_ ( .D(n9168), .CLK(clk), .Q(arr[866]) );
  DFFPOSX1 arr_reg_21__4_ ( .D(n9167), .CLK(clk), .Q(arr[865]) );
  DFFPOSX1 arr_reg_21__3_ ( .D(n9166), .CLK(clk), .Q(arr[864]) );
  DFFPOSX1 arr_reg_21__2_ ( .D(n9165), .CLK(clk), .Q(arr[863]) );
  DFFPOSX1 arr_reg_21__1_ ( .D(n9164), .CLK(clk), .Q(arr[862]) );
  DFFPOSX1 arr_reg_21__0_ ( .D(n9163), .CLK(clk), .Q(arr[861]) );
  DFFPOSX1 arr_reg_20__40_ ( .D(n9162), .CLK(clk), .Q(arr[860]) );
  DFFPOSX1 arr_reg_20__39_ ( .D(n9161), .CLK(clk), .Q(arr[859]) );
  DFFPOSX1 arr_reg_20__38_ ( .D(n9160), .CLK(clk), .Q(arr[858]) );
  DFFPOSX1 arr_reg_20__37_ ( .D(n9159), .CLK(clk), .Q(arr[857]) );
  DFFPOSX1 arr_reg_20__36_ ( .D(n9158), .CLK(clk), .Q(arr[856]) );
  DFFPOSX1 arr_reg_20__35_ ( .D(n9157), .CLK(clk), .Q(arr[855]) );
  DFFPOSX1 arr_reg_20__34_ ( .D(n9156), .CLK(clk), .Q(arr[854]) );
  DFFPOSX1 arr_reg_20__33_ ( .D(n9155), .CLK(clk), .Q(arr[853]) );
  DFFPOSX1 arr_reg_20__32_ ( .D(n9154), .CLK(clk), .Q(arr[852]) );
  DFFPOSX1 arr_reg_20__31_ ( .D(n9153), .CLK(clk), .Q(arr[851]) );
  DFFPOSX1 arr_reg_20__30_ ( .D(n9152), .CLK(clk), .Q(arr[850]) );
  DFFPOSX1 arr_reg_20__29_ ( .D(n9151), .CLK(clk), .Q(arr[849]) );
  DFFPOSX1 arr_reg_20__28_ ( .D(n9150), .CLK(clk), .Q(arr[848]) );
  DFFPOSX1 arr_reg_20__27_ ( .D(n9149), .CLK(clk), .Q(arr[847]) );
  DFFPOSX1 arr_reg_20__26_ ( .D(n9148), .CLK(clk), .Q(arr[846]) );
  DFFPOSX1 arr_reg_20__25_ ( .D(n9147), .CLK(clk), .Q(arr[845]) );
  DFFPOSX1 arr_reg_20__24_ ( .D(n9146), .CLK(clk), .Q(arr[844]) );
  DFFPOSX1 arr_reg_20__23_ ( .D(n9145), .CLK(clk), .Q(arr[843]) );
  DFFPOSX1 arr_reg_20__22_ ( .D(n9144), .CLK(clk), .Q(arr[842]) );
  DFFPOSX1 arr_reg_20__21_ ( .D(n9143), .CLK(clk), .Q(arr[841]) );
  DFFPOSX1 arr_reg_20__20_ ( .D(n9142), .CLK(clk), .Q(arr[840]) );
  DFFPOSX1 arr_reg_20__19_ ( .D(n9141), .CLK(clk), .Q(arr[839]) );
  DFFPOSX1 arr_reg_20__18_ ( .D(n9140), .CLK(clk), .Q(arr[838]) );
  DFFPOSX1 arr_reg_20__17_ ( .D(n9139), .CLK(clk), .Q(arr[837]) );
  DFFPOSX1 arr_reg_20__16_ ( .D(n9138), .CLK(clk), .Q(arr[836]) );
  DFFPOSX1 arr_reg_20__15_ ( .D(n9137), .CLK(clk), .Q(arr[835]) );
  DFFPOSX1 arr_reg_20__14_ ( .D(n9136), .CLK(clk), .Q(arr[834]) );
  DFFPOSX1 arr_reg_20__13_ ( .D(n9135), .CLK(clk), .Q(arr[833]) );
  DFFPOSX1 arr_reg_20__12_ ( .D(n9134), .CLK(clk), .Q(arr[832]) );
  DFFPOSX1 arr_reg_20__11_ ( .D(n9133), .CLK(clk), .Q(arr[831]) );
  DFFPOSX1 arr_reg_20__10_ ( .D(n9132), .CLK(clk), .Q(arr[830]) );
  DFFPOSX1 arr_reg_20__9_ ( .D(n9131), .CLK(clk), .Q(arr[829]) );
  DFFPOSX1 arr_reg_20__8_ ( .D(n9130), .CLK(clk), .Q(arr[828]) );
  DFFPOSX1 arr_reg_20__7_ ( .D(n9129), .CLK(clk), .Q(arr[827]) );
  DFFPOSX1 arr_reg_20__6_ ( .D(n9128), .CLK(clk), .Q(arr[826]) );
  DFFPOSX1 arr_reg_20__5_ ( .D(n9127), .CLK(clk), .Q(arr[825]) );
  DFFPOSX1 arr_reg_20__4_ ( .D(n9126), .CLK(clk), .Q(arr[824]) );
  DFFPOSX1 arr_reg_20__3_ ( .D(n9125), .CLK(clk), .Q(arr[823]) );
  DFFPOSX1 arr_reg_20__2_ ( .D(n9124), .CLK(clk), .Q(arr[822]) );
  DFFPOSX1 arr_reg_20__1_ ( .D(n9123), .CLK(clk), .Q(arr[821]) );
  DFFPOSX1 arr_reg_20__0_ ( .D(n9122), .CLK(clk), .Q(arr[820]) );
  DFFPOSX1 arr_reg_19__40_ ( .D(n9121), .CLK(clk), .Q(arr[819]) );
  DFFPOSX1 arr_reg_19__39_ ( .D(n9120), .CLK(clk), .Q(arr[818]) );
  DFFPOSX1 arr_reg_19__38_ ( .D(n9119), .CLK(clk), .Q(arr[817]) );
  DFFPOSX1 arr_reg_19__37_ ( .D(n9118), .CLK(clk), .Q(arr[816]) );
  DFFPOSX1 arr_reg_19__36_ ( .D(n9117), .CLK(clk), .Q(arr[815]) );
  DFFPOSX1 arr_reg_19__35_ ( .D(n9116), .CLK(clk), .Q(arr[814]) );
  DFFPOSX1 arr_reg_19__34_ ( .D(n9115), .CLK(clk), .Q(arr[813]) );
  DFFPOSX1 arr_reg_19__33_ ( .D(n9114), .CLK(clk), .Q(arr[812]) );
  DFFPOSX1 arr_reg_19__32_ ( .D(n9113), .CLK(clk), .Q(arr[811]) );
  DFFPOSX1 arr_reg_19__31_ ( .D(n9112), .CLK(clk), .Q(arr[810]) );
  DFFPOSX1 arr_reg_19__30_ ( .D(n9111), .CLK(clk), .Q(arr[809]) );
  DFFPOSX1 arr_reg_19__29_ ( .D(n9110), .CLK(clk), .Q(arr[808]) );
  DFFPOSX1 arr_reg_19__28_ ( .D(n9109), .CLK(clk), .Q(arr[807]) );
  DFFPOSX1 arr_reg_19__27_ ( .D(n9108), .CLK(clk), .Q(arr[806]) );
  DFFPOSX1 arr_reg_19__26_ ( .D(n9107), .CLK(clk), .Q(arr[805]) );
  DFFPOSX1 arr_reg_19__25_ ( .D(n9106), .CLK(clk), .Q(arr[804]) );
  DFFPOSX1 arr_reg_19__24_ ( .D(n9105), .CLK(clk), .Q(arr[803]) );
  DFFPOSX1 arr_reg_19__23_ ( .D(n9104), .CLK(clk), .Q(arr[802]) );
  DFFPOSX1 arr_reg_19__22_ ( .D(n9103), .CLK(clk), .Q(arr[801]) );
  DFFPOSX1 arr_reg_19__21_ ( .D(n9102), .CLK(clk), .Q(arr[800]) );
  DFFPOSX1 arr_reg_19__20_ ( .D(n9101), .CLK(clk), .Q(arr[799]) );
  DFFPOSX1 arr_reg_19__19_ ( .D(n9100), .CLK(clk), .Q(arr[798]) );
  DFFPOSX1 arr_reg_19__18_ ( .D(n9099), .CLK(clk), .Q(arr[797]) );
  DFFPOSX1 arr_reg_19__17_ ( .D(n9098), .CLK(clk), .Q(arr[796]) );
  DFFPOSX1 arr_reg_19__16_ ( .D(n9097), .CLK(clk), .Q(arr[795]) );
  DFFPOSX1 arr_reg_19__15_ ( .D(n9096), .CLK(clk), .Q(arr[794]) );
  DFFPOSX1 arr_reg_19__14_ ( .D(n9095), .CLK(clk), .Q(arr[793]) );
  DFFPOSX1 arr_reg_19__13_ ( .D(n9094), .CLK(clk), .Q(arr[792]) );
  DFFPOSX1 arr_reg_19__12_ ( .D(n9093), .CLK(clk), .Q(arr[791]) );
  DFFPOSX1 arr_reg_19__11_ ( .D(n9092), .CLK(clk), .Q(arr[790]) );
  DFFPOSX1 arr_reg_19__10_ ( .D(n9091), .CLK(clk), .Q(arr[789]) );
  DFFPOSX1 arr_reg_19__9_ ( .D(n9090), .CLK(clk), .Q(arr[788]) );
  DFFPOSX1 arr_reg_19__8_ ( .D(n9089), .CLK(clk), .Q(arr[787]) );
  DFFPOSX1 arr_reg_19__7_ ( .D(n9088), .CLK(clk), .Q(arr[786]) );
  DFFPOSX1 arr_reg_19__6_ ( .D(n9087), .CLK(clk), .Q(arr[785]) );
  DFFPOSX1 arr_reg_19__5_ ( .D(n9086), .CLK(clk), .Q(arr[784]) );
  DFFPOSX1 arr_reg_19__4_ ( .D(n9085), .CLK(clk), .Q(arr[783]) );
  DFFPOSX1 arr_reg_19__3_ ( .D(n9084), .CLK(clk), .Q(arr[782]) );
  DFFPOSX1 arr_reg_19__2_ ( .D(n9083), .CLK(clk), .Q(arr[781]) );
  DFFPOSX1 arr_reg_19__1_ ( .D(n9082), .CLK(clk), .Q(arr[780]) );
  DFFPOSX1 arr_reg_19__0_ ( .D(n9081), .CLK(clk), .Q(arr[779]) );
  DFFPOSX1 arr_reg_18__40_ ( .D(n9080), .CLK(clk), .Q(arr[778]) );
  DFFPOSX1 arr_reg_18__39_ ( .D(n9079), .CLK(clk), .Q(arr[777]) );
  DFFPOSX1 arr_reg_18__38_ ( .D(n9078), .CLK(clk), .Q(arr[776]) );
  DFFPOSX1 arr_reg_18__37_ ( .D(n9077), .CLK(clk), .Q(arr[775]) );
  DFFPOSX1 arr_reg_18__36_ ( .D(n9076), .CLK(clk), .Q(arr[774]) );
  DFFPOSX1 arr_reg_18__35_ ( .D(n9075), .CLK(clk), .Q(arr[773]) );
  DFFPOSX1 arr_reg_18__34_ ( .D(n9074), .CLK(clk), .Q(arr[772]) );
  DFFPOSX1 arr_reg_18__33_ ( .D(n9073), .CLK(clk), .Q(arr[771]) );
  DFFPOSX1 arr_reg_18__32_ ( .D(n9072), .CLK(clk), .Q(arr[770]) );
  DFFPOSX1 arr_reg_18__31_ ( .D(n9071), .CLK(clk), .Q(arr[769]) );
  DFFPOSX1 arr_reg_18__30_ ( .D(n9070), .CLK(clk), .Q(arr[768]) );
  DFFPOSX1 arr_reg_18__29_ ( .D(n9069), .CLK(clk), .Q(arr[767]) );
  DFFPOSX1 arr_reg_18__28_ ( .D(n9068), .CLK(clk), .Q(arr[766]) );
  DFFPOSX1 arr_reg_18__27_ ( .D(n9067), .CLK(clk), .Q(arr[765]) );
  DFFPOSX1 arr_reg_18__26_ ( .D(n9066), .CLK(clk), .Q(arr[764]) );
  DFFPOSX1 arr_reg_18__25_ ( .D(n9065), .CLK(clk), .Q(arr[763]) );
  DFFPOSX1 arr_reg_18__24_ ( .D(n9064), .CLK(clk), .Q(arr[762]) );
  DFFPOSX1 arr_reg_18__23_ ( .D(n9063), .CLK(clk), .Q(arr[761]) );
  DFFPOSX1 arr_reg_18__22_ ( .D(n9062), .CLK(clk), .Q(arr[760]) );
  DFFPOSX1 arr_reg_18__21_ ( .D(n9061), .CLK(clk), .Q(arr[759]) );
  DFFPOSX1 arr_reg_18__20_ ( .D(n9060), .CLK(clk), .Q(arr[758]) );
  DFFPOSX1 arr_reg_18__19_ ( .D(n9059), .CLK(clk), .Q(arr[757]) );
  DFFPOSX1 arr_reg_18__18_ ( .D(n9058), .CLK(clk), .Q(arr[756]) );
  DFFPOSX1 arr_reg_18__17_ ( .D(n9057), .CLK(clk), .Q(arr[755]) );
  DFFPOSX1 arr_reg_18__16_ ( .D(n9056), .CLK(clk), .Q(arr[754]) );
  DFFPOSX1 arr_reg_18__15_ ( .D(n9055), .CLK(clk), .Q(arr[753]) );
  DFFPOSX1 arr_reg_18__14_ ( .D(n9054), .CLK(clk), .Q(arr[752]) );
  DFFPOSX1 arr_reg_18__13_ ( .D(n9053), .CLK(clk), .Q(arr[751]) );
  DFFPOSX1 arr_reg_18__12_ ( .D(n9052), .CLK(clk), .Q(arr[750]) );
  DFFPOSX1 arr_reg_18__11_ ( .D(n9051), .CLK(clk), .Q(arr[749]) );
  DFFPOSX1 arr_reg_18__10_ ( .D(n9050), .CLK(clk), .Q(arr[748]) );
  DFFPOSX1 arr_reg_18__9_ ( .D(n9049), .CLK(clk), .Q(arr[747]) );
  DFFPOSX1 arr_reg_18__8_ ( .D(n9048), .CLK(clk), .Q(arr[746]) );
  DFFPOSX1 arr_reg_18__7_ ( .D(n9047), .CLK(clk), .Q(arr[745]) );
  DFFPOSX1 arr_reg_18__6_ ( .D(n9046), .CLK(clk), .Q(arr[744]) );
  DFFPOSX1 arr_reg_18__5_ ( .D(n9045), .CLK(clk), .Q(arr[743]) );
  DFFPOSX1 arr_reg_18__4_ ( .D(n9044), .CLK(clk), .Q(arr[742]) );
  DFFPOSX1 arr_reg_18__3_ ( .D(n9043), .CLK(clk), .Q(arr[741]) );
  DFFPOSX1 arr_reg_18__2_ ( .D(n9042), .CLK(clk), .Q(arr[740]) );
  DFFPOSX1 arr_reg_18__1_ ( .D(n9041), .CLK(clk), .Q(arr[739]) );
  DFFPOSX1 arr_reg_18__0_ ( .D(n9040), .CLK(clk), .Q(arr[738]) );
  DFFPOSX1 arr_reg_17__40_ ( .D(n9039), .CLK(clk), .Q(arr[737]) );
  DFFPOSX1 arr_reg_17__39_ ( .D(n9038), .CLK(clk), .Q(arr[736]) );
  DFFPOSX1 arr_reg_17__38_ ( .D(n9037), .CLK(clk), .Q(arr[735]) );
  DFFPOSX1 arr_reg_17__37_ ( .D(n9036), .CLK(clk), .Q(arr[734]) );
  DFFPOSX1 arr_reg_17__36_ ( .D(n9035), .CLK(clk), .Q(arr[733]) );
  DFFPOSX1 arr_reg_17__35_ ( .D(n9034), .CLK(clk), .Q(arr[732]) );
  DFFPOSX1 arr_reg_17__34_ ( .D(n9033), .CLK(clk), .Q(arr[731]) );
  DFFPOSX1 arr_reg_17__33_ ( .D(n9032), .CLK(clk), .Q(arr[730]) );
  DFFPOSX1 arr_reg_17__32_ ( .D(n9031), .CLK(clk), .Q(arr[729]) );
  DFFPOSX1 arr_reg_17__31_ ( .D(n9030), .CLK(clk), .Q(arr[728]) );
  DFFPOSX1 arr_reg_17__30_ ( .D(n9029), .CLK(clk), .Q(arr[727]) );
  DFFPOSX1 arr_reg_17__29_ ( .D(n9028), .CLK(clk), .Q(arr[726]) );
  DFFPOSX1 arr_reg_17__28_ ( .D(n9027), .CLK(clk), .Q(arr[725]) );
  DFFPOSX1 arr_reg_17__27_ ( .D(n9026), .CLK(clk), .Q(arr[724]) );
  DFFPOSX1 arr_reg_17__26_ ( .D(n9025), .CLK(clk), .Q(arr[723]) );
  DFFPOSX1 arr_reg_17__25_ ( .D(n9024), .CLK(clk), .Q(arr[722]) );
  DFFPOSX1 arr_reg_17__24_ ( .D(n9023), .CLK(clk), .Q(arr[721]) );
  DFFPOSX1 arr_reg_17__23_ ( .D(n9022), .CLK(clk), .Q(arr[720]) );
  DFFPOSX1 arr_reg_17__22_ ( .D(n9021), .CLK(clk), .Q(arr[719]) );
  DFFPOSX1 arr_reg_17__21_ ( .D(n9020), .CLK(clk), .Q(arr[718]) );
  DFFPOSX1 arr_reg_17__20_ ( .D(n9019), .CLK(clk), .Q(arr[717]) );
  DFFPOSX1 arr_reg_17__19_ ( .D(n9018), .CLK(clk), .Q(arr[716]) );
  DFFPOSX1 arr_reg_17__18_ ( .D(n9017), .CLK(clk), .Q(arr[715]) );
  DFFPOSX1 arr_reg_17__17_ ( .D(n9016), .CLK(clk), .Q(arr[714]) );
  DFFPOSX1 arr_reg_17__16_ ( .D(n9015), .CLK(clk), .Q(arr[713]) );
  DFFPOSX1 arr_reg_17__15_ ( .D(n9014), .CLK(clk), .Q(arr[712]) );
  DFFPOSX1 arr_reg_17__14_ ( .D(n9013), .CLK(clk), .Q(arr[711]) );
  DFFPOSX1 arr_reg_17__13_ ( .D(n9012), .CLK(clk), .Q(arr[710]) );
  DFFPOSX1 arr_reg_17__12_ ( .D(n9011), .CLK(clk), .Q(arr[709]) );
  DFFPOSX1 arr_reg_17__11_ ( .D(n9010), .CLK(clk), .Q(arr[708]) );
  DFFPOSX1 arr_reg_17__10_ ( .D(n9009), .CLK(clk), .Q(arr[707]) );
  DFFPOSX1 arr_reg_17__9_ ( .D(n9008), .CLK(clk), .Q(arr[706]) );
  DFFPOSX1 arr_reg_17__8_ ( .D(n9007), .CLK(clk), .Q(arr[705]) );
  DFFPOSX1 arr_reg_17__7_ ( .D(n9006), .CLK(clk), .Q(arr[704]) );
  DFFPOSX1 arr_reg_17__6_ ( .D(n9005), .CLK(clk), .Q(arr[703]) );
  DFFPOSX1 arr_reg_17__5_ ( .D(n9004), .CLK(clk), .Q(arr[702]) );
  DFFPOSX1 arr_reg_17__4_ ( .D(n9003), .CLK(clk), .Q(arr[701]) );
  DFFPOSX1 arr_reg_17__3_ ( .D(n9002), .CLK(clk), .Q(arr[700]) );
  DFFPOSX1 arr_reg_17__2_ ( .D(n9001), .CLK(clk), .Q(arr[699]) );
  DFFPOSX1 arr_reg_17__1_ ( .D(n9000), .CLK(clk), .Q(arr[698]) );
  DFFPOSX1 arr_reg_17__0_ ( .D(n8999), .CLK(clk), .Q(arr[697]) );
  DFFPOSX1 arr_reg_16__40_ ( .D(n8998), .CLK(clk), .Q(arr[696]) );
  DFFPOSX1 arr_reg_16__39_ ( .D(n8997), .CLK(clk), .Q(arr[695]) );
  DFFPOSX1 arr_reg_16__38_ ( .D(n8996), .CLK(clk), .Q(arr[694]) );
  DFFPOSX1 arr_reg_16__37_ ( .D(n8995), .CLK(clk), .Q(arr[693]) );
  DFFPOSX1 arr_reg_16__36_ ( .D(n8994), .CLK(clk), .Q(arr[692]) );
  DFFPOSX1 arr_reg_16__35_ ( .D(n8993), .CLK(clk), .Q(arr[691]) );
  DFFPOSX1 arr_reg_16__34_ ( .D(n8992), .CLK(clk), .Q(arr[690]) );
  DFFPOSX1 arr_reg_16__33_ ( .D(n8991), .CLK(clk), .Q(arr[689]) );
  DFFPOSX1 arr_reg_16__32_ ( .D(n8990), .CLK(clk), .Q(arr[688]) );
  DFFPOSX1 arr_reg_16__31_ ( .D(n8989), .CLK(clk), .Q(arr[687]) );
  DFFPOSX1 arr_reg_16__30_ ( .D(n8988), .CLK(clk), .Q(arr[686]) );
  DFFPOSX1 arr_reg_16__29_ ( .D(n8987), .CLK(clk), .Q(arr[685]) );
  DFFPOSX1 arr_reg_16__28_ ( .D(n8986), .CLK(clk), .Q(arr[684]) );
  DFFPOSX1 arr_reg_16__27_ ( .D(n8985), .CLK(clk), .Q(arr[683]) );
  DFFPOSX1 arr_reg_16__26_ ( .D(n8984), .CLK(clk), .Q(arr[682]) );
  DFFPOSX1 arr_reg_16__25_ ( .D(n8983), .CLK(clk), .Q(arr[681]) );
  DFFPOSX1 arr_reg_16__24_ ( .D(n8982), .CLK(clk), .Q(arr[680]) );
  DFFPOSX1 arr_reg_16__23_ ( .D(n8981), .CLK(clk), .Q(arr[679]) );
  DFFPOSX1 arr_reg_16__22_ ( .D(n8980), .CLK(clk), .Q(arr[678]) );
  DFFPOSX1 arr_reg_16__21_ ( .D(n8979), .CLK(clk), .Q(arr[677]) );
  DFFPOSX1 arr_reg_16__20_ ( .D(n8978), .CLK(clk), .Q(arr[676]) );
  DFFPOSX1 arr_reg_16__19_ ( .D(n8977), .CLK(clk), .Q(arr[675]) );
  DFFPOSX1 arr_reg_16__18_ ( .D(n8976), .CLK(clk), .Q(arr[674]) );
  DFFPOSX1 arr_reg_16__17_ ( .D(n8975), .CLK(clk), .Q(arr[673]) );
  DFFPOSX1 arr_reg_16__16_ ( .D(n8974), .CLK(clk), .Q(arr[672]) );
  DFFPOSX1 arr_reg_16__15_ ( .D(n8973), .CLK(clk), .Q(arr[671]) );
  DFFPOSX1 arr_reg_16__14_ ( .D(n8972), .CLK(clk), .Q(arr[670]) );
  DFFPOSX1 arr_reg_16__13_ ( .D(n8971), .CLK(clk), .Q(arr[669]) );
  DFFPOSX1 arr_reg_16__12_ ( .D(n8970), .CLK(clk), .Q(arr[668]) );
  DFFPOSX1 arr_reg_16__11_ ( .D(n8969), .CLK(clk), .Q(arr[667]) );
  DFFPOSX1 arr_reg_16__10_ ( .D(n8968), .CLK(clk), .Q(arr[666]) );
  DFFPOSX1 arr_reg_16__9_ ( .D(n8967), .CLK(clk), .Q(arr[665]) );
  DFFPOSX1 arr_reg_16__8_ ( .D(n8966), .CLK(clk), .Q(arr[664]) );
  DFFPOSX1 arr_reg_16__7_ ( .D(n8965), .CLK(clk), .Q(arr[663]) );
  DFFPOSX1 arr_reg_16__6_ ( .D(n8964), .CLK(clk), .Q(arr[662]) );
  DFFPOSX1 arr_reg_16__5_ ( .D(n8963), .CLK(clk), .Q(arr[661]) );
  DFFPOSX1 arr_reg_16__4_ ( .D(n8962), .CLK(clk), .Q(arr[660]) );
  DFFPOSX1 arr_reg_16__3_ ( .D(n8961), .CLK(clk), .Q(arr[659]) );
  DFFPOSX1 arr_reg_16__2_ ( .D(n8960), .CLK(clk), .Q(arr[658]) );
  DFFPOSX1 arr_reg_16__1_ ( .D(n8959), .CLK(clk), .Q(arr[657]) );
  DFFPOSX1 arr_reg_16__0_ ( .D(n8958), .CLK(clk), .Q(arr[656]) );
  DFFPOSX1 arr_reg_15__40_ ( .D(n8957), .CLK(clk), .Q(arr[655]) );
  DFFPOSX1 arr_reg_15__39_ ( .D(n8956), .CLK(clk), .Q(arr[654]) );
  DFFPOSX1 arr_reg_15__38_ ( .D(n8955), .CLK(clk), .Q(arr[653]) );
  DFFPOSX1 arr_reg_15__37_ ( .D(n8954), .CLK(clk), .Q(arr[652]) );
  DFFPOSX1 arr_reg_15__36_ ( .D(n8953), .CLK(clk), .Q(arr[651]) );
  DFFPOSX1 arr_reg_15__35_ ( .D(n8952), .CLK(clk), .Q(arr[650]) );
  DFFPOSX1 arr_reg_15__34_ ( .D(n8951), .CLK(clk), .Q(arr[649]) );
  DFFPOSX1 arr_reg_15__33_ ( .D(n8950), .CLK(clk), .Q(arr[648]) );
  DFFPOSX1 arr_reg_15__32_ ( .D(n8949), .CLK(clk), .Q(arr[647]) );
  DFFPOSX1 arr_reg_15__31_ ( .D(n8948), .CLK(clk), .Q(arr[646]) );
  DFFPOSX1 arr_reg_15__30_ ( .D(n8947), .CLK(clk), .Q(arr[645]) );
  DFFPOSX1 arr_reg_15__29_ ( .D(n8946), .CLK(clk), .Q(arr[644]) );
  DFFPOSX1 arr_reg_15__28_ ( .D(n8945), .CLK(clk), .Q(arr[643]) );
  DFFPOSX1 arr_reg_15__27_ ( .D(n8944), .CLK(clk), .Q(arr[642]) );
  DFFPOSX1 arr_reg_15__26_ ( .D(n8943), .CLK(clk), .Q(arr[641]) );
  DFFPOSX1 arr_reg_15__25_ ( .D(n8942), .CLK(clk), .Q(arr[640]) );
  DFFPOSX1 arr_reg_15__24_ ( .D(n8941), .CLK(clk), .Q(arr[639]) );
  DFFPOSX1 arr_reg_15__23_ ( .D(n8940), .CLK(clk), .Q(arr[638]) );
  DFFPOSX1 arr_reg_15__22_ ( .D(n8939), .CLK(clk), .Q(arr[637]) );
  DFFPOSX1 arr_reg_15__21_ ( .D(n8938), .CLK(clk), .Q(arr[636]) );
  DFFPOSX1 arr_reg_15__20_ ( .D(n8937), .CLK(clk), .Q(arr[635]) );
  DFFPOSX1 arr_reg_15__19_ ( .D(n8936), .CLK(clk), .Q(arr[634]) );
  DFFPOSX1 arr_reg_15__18_ ( .D(n8935), .CLK(clk), .Q(arr[633]) );
  DFFPOSX1 arr_reg_15__17_ ( .D(n8934), .CLK(clk), .Q(arr[632]) );
  DFFPOSX1 arr_reg_15__16_ ( .D(n8933), .CLK(clk), .Q(arr[631]) );
  DFFPOSX1 arr_reg_15__15_ ( .D(n8932), .CLK(clk), .Q(arr[630]) );
  DFFPOSX1 arr_reg_15__14_ ( .D(n8931), .CLK(clk), .Q(arr[629]) );
  DFFPOSX1 arr_reg_15__13_ ( .D(n8930), .CLK(clk), .Q(arr[628]) );
  DFFPOSX1 arr_reg_15__12_ ( .D(n8929), .CLK(clk), .Q(arr[627]) );
  DFFPOSX1 arr_reg_15__11_ ( .D(n8928), .CLK(clk), .Q(arr[626]) );
  DFFPOSX1 arr_reg_15__10_ ( .D(n8927), .CLK(clk), .Q(arr[625]) );
  DFFPOSX1 arr_reg_15__9_ ( .D(n8926), .CLK(clk), .Q(arr[624]) );
  DFFPOSX1 arr_reg_15__8_ ( .D(n8925), .CLK(clk), .Q(arr[623]) );
  DFFPOSX1 arr_reg_15__7_ ( .D(n8924), .CLK(clk), .Q(arr[622]) );
  DFFPOSX1 arr_reg_15__6_ ( .D(n8923), .CLK(clk), .Q(arr[621]) );
  DFFPOSX1 arr_reg_15__5_ ( .D(n8922), .CLK(clk), .Q(arr[620]) );
  DFFPOSX1 arr_reg_15__4_ ( .D(n8921), .CLK(clk), .Q(arr[619]) );
  DFFPOSX1 arr_reg_15__3_ ( .D(n8920), .CLK(clk), .Q(arr[618]) );
  DFFPOSX1 arr_reg_15__2_ ( .D(n8919), .CLK(clk), .Q(arr[617]) );
  DFFPOSX1 arr_reg_15__1_ ( .D(n8918), .CLK(clk), .Q(arr[616]) );
  DFFPOSX1 arr_reg_15__0_ ( .D(n8917), .CLK(clk), .Q(arr[615]) );
  DFFPOSX1 arr_reg_14__40_ ( .D(n8916), .CLK(clk), .Q(arr[614]) );
  DFFPOSX1 arr_reg_14__39_ ( .D(n8915), .CLK(clk), .Q(arr[613]) );
  DFFPOSX1 arr_reg_14__38_ ( .D(n8914), .CLK(clk), .Q(arr[612]) );
  DFFPOSX1 arr_reg_14__37_ ( .D(n8913), .CLK(clk), .Q(arr[611]) );
  DFFPOSX1 arr_reg_14__36_ ( .D(n8912), .CLK(clk), .Q(arr[610]) );
  DFFPOSX1 arr_reg_14__35_ ( .D(n8911), .CLK(clk), .Q(arr[609]) );
  DFFPOSX1 arr_reg_14__34_ ( .D(n8910), .CLK(clk), .Q(arr[608]) );
  DFFPOSX1 arr_reg_14__33_ ( .D(n8909), .CLK(clk), .Q(arr[607]) );
  DFFPOSX1 arr_reg_14__32_ ( .D(n8908), .CLK(clk), .Q(arr[606]) );
  DFFPOSX1 arr_reg_14__31_ ( .D(n8907), .CLK(clk), .Q(arr[605]) );
  DFFPOSX1 arr_reg_14__30_ ( .D(n8906), .CLK(clk), .Q(arr[604]) );
  DFFPOSX1 arr_reg_14__29_ ( .D(n8905), .CLK(clk), .Q(arr[603]) );
  DFFPOSX1 arr_reg_14__28_ ( .D(n8904), .CLK(clk), .Q(arr[602]) );
  DFFPOSX1 arr_reg_14__27_ ( .D(n8903), .CLK(clk), .Q(arr[601]) );
  DFFPOSX1 arr_reg_14__26_ ( .D(n8902), .CLK(clk), .Q(arr[600]) );
  DFFPOSX1 arr_reg_14__25_ ( .D(n8901), .CLK(clk), .Q(arr[599]) );
  DFFPOSX1 arr_reg_14__24_ ( .D(n8900), .CLK(clk), .Q(arr[598]) );
  DFFPOSX1 arr_reg_14__23_ ( .D(n8899), .CLK(clk), .Q(arr[597]) );
  DFFPOSX1 arr_reg_14__22_ ( .D(n8898), .CLK(clk), .Q(arr[596]) );
  DFFPOSX1 arr_reg_14__21_ ( .D(n8897), .CLK(clk), .Q(arr[595]) );
  DFFPOSX1 arr_reg_14__20_ ( .D(n8896), .CLK(clk), .Q(arr[594]) );
  DFFPOSX1 arr_reg_14__19_ ( .D(n8895), .CLK(clk), .Q(arr[593]) );
  DFFPOSX1 arr_reg_14__18_ ( .D(n8894), .CLK(clk), .Q(arr[592]) );
  DFFPOSX1 arr_reg_14__17_ ( .D(n8893), .CLK(clk), .Q(arr[591]) );
  DFFPOSX1 arr_reg_14__16_ ( .D(n8892), .CLK(clk), .Q(arr[590]) );
  DFFPOSX1 arr_reg_14__15_ ( .D(n8891), .CLK(clk), .Q(arr[589]) );
  DFFPOSX1 arr_reg_14__14_ ( .D(n8890), .CLK(clk), .Q(arr[588]) );
  DFFPOSX1 arr_reg_14__13_ ( .D(n8889), .CLK(clk), .Q(arr[587]) );
  DFFPOSX1 arr_reg_14__12_ ( .D(n8888), .CLK(clk), .Q(arr[586]) );
  DFFPOSX1 arr_reg_14__11_ ( .D(n8887), .CLK(clk), .Q(arr[585]) );
  DFFPOSX1 arr_reg_14__10_ ( .D(n8886), .CLK(clk), .Q(arr[584]) );
  DFFPOSX1 arr_reg_14__9_ ( .D(n8885), .CLK(clk), .Q(arr[583]) );
  DFFPOSX1 arr_reg_14__8_ ( .D(n8884), .CLK(clk), .Q(arr[582]) );
  DFFPOSX1 arr_reg_14__7_ ( .D(n8883), .CLK(clk), .Q(arr[581]) );
  DFFPOSX1 arr_reg_14__6_ ( .D(n8882), .CLK(clk), .Q(arr[580]) );
  DFFPOSX1 arr_reg_14__5_ ( .D(n8881), .CLK(clk), .Q(arr[579]) );
  DFFPOSX1 arr_reg_14__4_ ( .D(n8880), .CLK(clk), .Q(arr[578]) );
  DFFPOSX1 arr_reg_14__3_ ( .D(n8879), .CLK(clk), .Q(arr[577]) );
  DFFPOSX1 arr_reg_14__2_ ( .D(n8878), .CLK(clk), .Q(arr[576]) );
  DFFPOSX1 arr_reg_14__1_ ( .D(n8877), .CLK(clk), .Q(arr[575]) );
  DFFPOSX1 arr_reg_14__0_ ( .D(n8876), .CLK(clk), .Q(arr[574]) );
  DFFPOSX1 arr_reg_13__40_ ( .D(n8875), .CLK(clk), .Q(arr[573]) );
  DFFPOSX1 arr_reg_13__39_ ( .D(n8874), .CLK(clk), .Q(arr[572]) );
  DFFPOSX1 arr_reg_13__38_ ( .D(n8873), .CLK(clk), .Q(arr[571]) );
  DFFPOSX1 arr_reg_13__37_ ( .D(n8872), .CLK(clk), .Q(arr[570]) );
  DFFPOSX1 arr_reg_13__36_ ( .D(n8871), .CLK(clk), .Q(arr[569]) );
  DFFPOSX1 arr_reg_13__35_ ( .D(n8870), .CLK(clk), .Q(arr[568]) );
  DFFPOSX1 arr_reg_13__34_ ( .D(n8869), .CLK(clk), .Q(arr[567]) );
  DFFPOSX1 arr_reg_13__33_ ( .D(n8868), .CLK(clk), .Q(arr[566]) );
  DFFPOSX1 arr_reg_13__32_ ( .D(n8867), .CLK(clk), .Q(arr[565]) );
  DFFPOSX1 arr_reg_13__31_ ( .D(n8866), .CLK(clk), .Q(arr[564]) );
  DFFPOSX1 arr_reg_13__30_ ( .D(n8865), .CLK(clk), .Q(arr[563]) );
  DFFPOSX1 arr_reg_13__29_ ( .D(n8864), .CLK(clk), .Q(arr[562]) );
  DFFPOSX1 arr_reg_13__28_ ( .D(n8863), .CLK(clk), .Q(arr[561]) );
  DFFPOSX1 arr_reg_13__27_ ( .D(n8862), .CLK(clk), .Q(arr[560]) );
  DFFPOSX1 arr_reg_13__26_ ( .D(n8861), .CLK(clk), .Q(arr[559]) );
  DFFPOSX1 arr_reg_13__25_ ( .D(n8860), .CLK(clk), .Q(arr[558]) );
  DFFPOSX1 arr_reg_13__24_ ( .D(n8859), .CLK(clk), .Q(arr[557]) );
  DFFPOSX1 arr_reg_13__23_ ( .D(n8858), .CLK(clk), .Q(arr[556]) );
  DFFPOSX1 arr_reg_13__22_ ( .D(n8857), .CLK(clk), .Q(arr[555]) );
  DFFPOSX1 arr_reg_13__21_ ( .D(n8856), .CLK(clk), .Q(arr[554]) );
  DFFPOSX1 arr_reg_13__20_ ( .D(n8855), .CLK(clk), .Q(arr[553]) );
  DFFPOSX1 arr_reg_13__19_ ( .D(n8854), .CLK(clk), .Q(arr[552]) );
  DFFPOSX1 arr_reg_13__18_ ( .D(n8853), .CLK(clk), .Q(arr[551]) );
  DFFPOSX1 arr_reg_13__17_ ( .D(n8852), .CLK(clk), .Q(arr[550]) );
  DFFPOSX1 arr_reg_13__16_ ( .D(n8851), .CLK(clk), .Q(arr[549]) );
  DFFPOSX1 arr_reg_13__15_ ( .D(n8850), .CLK(clk), .Q(arr[548]) );
  DFFPOSX1 arr_reg_13__14_ ( .D(n8849), .CLK(clk), .Q(arr[547]) );
  DFFPOSX1 arr_reg_13__13_ ( .D(n8848), .CLK(clk), .Q(arr[546]) );
  DFFPOSX1 arr_reg_13__12_ ( .D(n8847), .CLK(clk), .Q(arr[545]) );
  DFFPOSX1 arr_reg_13__11_ ( .D(n8846), .CLK(clk), .Q(arr[544]) );
  DFFPOSX1 arr_reg_13__10_ ( .D(n8845), .CLK(clk), .Q(arr[543]) );
  DFFPOSX1 arr_reg_13__9_ ( .D(n8844), .CLK(clk), .Q(arr[542]) );
  DFFPOSX1 arr_reg_13__8_ ( .D(n8843), .CLK(clk), .Q(arr[541]) );
  DFFPOSX1 arr_reg_13__7_ ( .D(n8842), .CLK(clk), .Q(arr[540]) );
  DFFPOSX1 arr_reg_13__6_ ( .D(n8841), .CLK(clk), .Q(arr[539]) );
  DFFPOSX1 arr_reg_13__5_ ( .D(n8840), .CLK(clk), .Q(arr[538]) );
  DFFPOSX1 arr_reg_13__4_ ( .D(n8839), .CLK(clk), .Q(arr[537]) );
  DFFPOSX1 arr_reg_13__3_ ( .D(n8838), .CLK(clk), .Q(arr[536]) );
  DFFPOSX1 arr_reg_13__2_ ( .D(n8837), .CLK(clk), .Q(arr[535]) );
  DFFPOSX1 arr_reg_13__1_ ( .D(n8836), .CLK(clk), .Q(arr[534]) );
  DFFPOSX1 arr_reg_13__0_ ( .D(n8835), .CLK(clk), .Q(arr[533]) );
  DFFPOSX1 arr_reg_12__40_ ( .D(n8834), .CLK(clk), .Q(arr[532]) );
  DFFPOSX1 arr_reg_12__39_ ( .D(n8833), .CLK(clk), .Q(arr[531]) );
  DFFPOSX1 arr_reg_12__38_ ( .D(n8832), .CLK(clk), .Q(arr[530]) );
  DFFPOSX1 arr_reg_12__37_ ( .D(n8831), .CLK(clk), .Q(arr[529]) );
  DFFPOSX1 arr_reg_12__36_ ( .D(n8830), .CLK(clk), .Q(arr[528]) );
  DFFPOSX1 arr_reg_12__35_ ( .D(n8829), .CLK(clk), .Q(arr[527]) );
  DFFPOSX1 arr_reg_12__34_ ( .D(n8828), .CLK(clk), .Q(arr[526]) );
  DFFPOSX1 arr_reg_12__33_ ( .D(n8827), .CLK(clk), .Q(arr[525]) );
  DFFPOSX1 arr_reg_12__32_ ( .D(n8826), .CLK(clk), .Q(arr[524]) );
  DFFPOSX1 arr_reg_12__31_ ( .D(n8825), .CLK(clk), .Q(arr[523]) );
  DFFPOSX1 arr_reg_12__30_ ( .D(n8824), .CLK(clk), .Q(arr[522]) );
  DFFPOSX1 arr_reg_12__29_ ( .D(n8823), .CLK(clk), .Q(arr[521]) );
  DFFPOSX1 arr_reg_12__28_ ( .D(n8822), .CLK(clk), .Q(arr[520]) );
  DFFPOSX1 arr_reg_12__27_ ( .D(n8821), .CLK(clk), .Q(arr[519]) );
  DFFPOSX1 arr_reg_12__26_ ( .D(n8820), .CLK(clk), .Q(arr[518]) );
  DFFPOSX1 arr_reg_12__25_ ( .D(n8819), .CLK(clk), .Q(arr[517]) );
  DFFPOSX1 arr_reg_12__24_ ( .D(n8818), .CLK(clk), .Q(arr[516]) );
  DFFPOSX1 arr_reg_12__23_ ( .D(n8817), .CLK(clk), .Q(arr[515]) );
  DFFPOSX1 arr_reg_12__22_ ( .D(n8816), .CLK(clk), .Q(arr[514]) );
  DFFPOSX1 arr_reg_12__21_ ( .D(n8815), .CLK(clk), .Q(arr[513]) );
  DFFPOSX1 arr_reg_12__20_ ( .D(n8814), .CLK(clk), .Q(arr[512]) );
  DFFPOSX1 arr_reg_12__19_ ( .D(n8813), .CLK(clk), .Q(arr[511]) );
  DFFPOSX1 arr_reg_12__18_ ( .D(n8812), .CLK(clk), .Q(arr[510]) );
  DFFPOSX1 arr_reg_12__17_ ( .D(n8811), .CLK(clk), .Q(arr[509]) );
  DFFPOSX1 arr_reg_12__16_ ( .D(n8810), .CLK(clk), .Q(arr[508]) );
  DFFPOSX1 arr_reg_12__15_ ( .D(n8809), .CLK(clk), .Q(arr[507]) );
  DFFPOSX1 arr_reg_12__14_ ( .D(n8808), .CLK(clk), .Q(arr[506]) );
  DFFPOSX1 arr_reg_12__13_ ( .D(n8807), .CLK(clk), .Q(arr[505]) );
  DFFPOSX1 arr_reg_12__12_ ( .D(n8806), .CLK(clk), .Q(arr[504]) );
  DFFPOSX1 arr_reg_12__11_ ( .D(n8805), .CLK(clk), .Q(arr[503]) );
  DFFPOSX1 arr_reg_12__10_ ( .D(n8804), .CLK(clk), .Q(arr[502]) );
  DFFPOSX1 arr_reg_12__9_ ( .D(n8803), .CLK(clk), .Q(arr[501]) );
  DFFPOSX1 arr_reg_12__8_ ( .D(n8802), .CLK(clk), .Q(arr[500]) );
  DFFPOSX1 arr_reg_12__7_ ( .D(n8801), .CLK(clk), .Q(arr[499]) );
  DFFPOSX1 arr_reg_12__6_ ( .D(n8800), .CLK(clk), .Q(arr[498]) );
  DFFPOSX1 arr_reg_12__5_ ( .D(n8799), .CLK(clk), .Q(arr[497]) );
  DFFPOSX1 arr_reg_12__4_ ( .D(n8798), .CLK(clk), .Q(arr[496]) );
  DFFPOSX1 arr_reg_12__3_ ( .D(n8797), .CLK(clk), .Q(arr[495]) );
  DFFPOSX1 arr_reg_12__2_ ( .D(n8796), .CLK(clk), .Q(arr[494]) );
  DFFPOSX1 arr_reg_12__1_ ( .D(n8795), .CLK(clk), .Q(arr[493]) );
  DFFPOSX1 arr_reg_12__0_ ( .D(n8794), .CLK(clk), .Q(arr[492]) );
  DFFPOSX1 arr_reg_11__40_ ( .D(n8793), .CLK(clk), .Q(arr[491]) );
  DFFPOSX1 arr_reg_11__39_ ( .D(n8792), .CLK(clk), .Q(arr[490]) );
  DFFPOSX1 arr_reg_11__38_ ( .D(n8791), .CLK(clk), .Q(arr[489]) );
  DFFPOSX1 arr_reg_11__37_ ( .D(n8790), .CLK(clk), .Q(arr[488]) );
  DFFPOSX1 arr_reg_11__36_ ( .D(n8789), .CLK(clk), .Q(arr[487]) );
  DFFPOSX1 arr_reg_11__35_ ( .D(n8788), .CLK(clk), .Q(arr[486]) );
  DFFPOSX1 arr_reg_11__34_ ( .D(n8787), .CLK(clk), .Q(arr[485]) );
  DFFPOSX1 arr_reg_11__33_ ( .D(n8786), .CLK(clk), .Q(arr[484]) );
  DFFPOSX1 arr_reg_11__32_ ( .D(n8785), .CLK(clk), .Q(arr[483]) );
  DFFPOSX1 arr_reg_11__31_ ( .D(n8784), .CLK(clk), .Q(arr[482]) );
  DFFPOSX1 arr_reg_11__30_ ( .D(n8783), .CLK(clk), .Q(arr[481]) );
  DFFPOSX1 arr_reg_11__29_ ( .D(n8782), .CLK(clk), .Q(arr[480]) );
  DFFPOSX1 arr_reg_11__28_ ( .D(n8781), .CLK(clk), .Q(arr[479]) );
  DFFPOSX1 arr_reg_11__27_ ( .D(n8780), .CLK(clk), .Q(arr[478]) );
  DFFPOSX1 arr_reg_11__26_ ( .D(n8779), .CLK(clk), .Q(arr[477]) );
  DFFPOSX1 arr_reg_11__25_ ( .D(n8778), .CLK(clk), .Q(arr[476]) );
  DFFPOSX1 arr_reg_11__24_ ( .D(n8777), .CLK(clk), .Q(arr[475]) );
  DFFPOSX1 arr_reg_11__23_ ( .D(n8776), .CLK(clk), .Q(arr[474]) );
  DFFPOSX1 arr_reg_11__22_ ( .D(n8775), .CLK(clk), .Q(arr[473]) );
  DFFPOSX1 arr_reg_11__21_ ( .D(n8774), .CLK(clk), .Q(arr[472]) );
  DFFPOSX1 arr_reg_11__20_ ( .D(n8773), .CLK(clk), .Q(arr[471]) );
  DFFPOSX1 arr_reg_11__19_ ( .D(n8772), .CLK(clk), .Q(arr[470]) );
  DFFPOSX1 arr_reg_11__18_ ( .D(n8771), .CLK(clk), .Q(arr[469]) );
  DFFPOSX1 arr_reg_11__17_ ( .D(n8770), .CLK(clk), .Q(arr[468]) );
  DFFPOSX1 arr_reg_11__16_ ( .D(n8769), .CLK(clk), .Q(arr[467]) );
  DFFPOSX1 arr_reg_11__15_ ( .D(n8768), .CLK(clk), .Q(arr[466]) );
  DFFPOSX1 arr_reg_11__14_ ( .D(n8767), .CLK(clk), .Q(arr[465]) );
  DFFPOSX1 arr_reg_11__13_ ( .D(n8766), .CLK(clk), .Q(arr[464]) );
  DFFPOSX1 arr_reg_11__12_ ( .D(n8765), .CLK(clk), .Q(arr[463]) );
  DFFPOSX1 arr_reg_11__11_ ( .D(n8764), .CLK(clk), .Q(arr[462]) );
  DFFPOSX1 arr_reg_11__10_ ( .D(n8763), .CLK(clk), .Q(arr[461]) );
  DFFPOSX1 arr_reg_11__9_ ( .D(n8762), .CLK(clk), .Q(arr[460]) );
  DFFPOSX1 arr_reg_11__8_ ( .D(n8761), .CLK(clk), .Q(arr[459]) );
  DFFPOSX1 arr_reg_11__7_ ( .D(n8760), .CLK(clk), .Q(arr[458]) );
  DFFPOSX1 arr_reg_11__6_ ( .D(n8759), .CLK(clk), .Q(arr[457]) );
  DFFPOSX1 arr_reg_11__5_ ( .D(n8758), .CLK(clk), .Q(arr[456]) );
  DFFPOSX1 arr_reg_11__4_ ( .D(n8757), .CLK(clk), .Q(arr[455]) );
  DFFPOSX1 arr_reg_11__3_ ( .D(n8756), .CLK(clk), .Q(arr[454]) );
  DFFPOSX1 arr_reg_11__2_ ( .D(n8755), .CLK(clk), .Q(arr[453]) );
  DFFPOSX1 arr_reg_11__1_ ( .D(n8754), .CLK(clk), .Q(arr[452]) );
  DFFPOSX1 arr_reg_11__0_ ( .D(n8753), .CLK(clk), .Q(arr[451]) );
  DFFPOSX1 arr_reg_10__40_ ( .D(n8752), .CLK(clk), .Q(arr[450]) );
  DFFPOSX1 arr_reg_10__39_ ( .D(n8751), .CLK(clk), .Q(arr[449]) );
  DFFPOSX1 arr_reg_10__38_ ( .D(n8750), .CLK(clk), .Q(arr[448]) );
  DFFPOSX1 arr_reg_10__37_ ( .D(n8749), .CLK(clk), .Q(arr[447]) );
  DFFPOSX1 arr_reg_10__36_ ( .D(n8748), .CLK(clk), .Q(arr[446]) );
  DFFPOSX1 arr_reg_10__35_ ( .D(n8747), .CLK(clk), .Q(arr[445]) );
  DFFPOSX1 arr_reg_10__34_ ( .D(n8746), .CLK(clk), .Q(arr[444]) );
  DFFPOSX1 arr_reg_10__33_ ( .D(n8745), .CLK(clk), .Q(arr[443]) );
  DFFPOSX1 arr_reg_10__32_ ( .D(n8744), .CLK(clk), .Q(arr[442]) );
  DFFPOSX1 arr_reg_10__31_ ( .D(n8743), .CLK(clk), .Q(arr[441]) );
  DFFPOSX1 arr_reg_10__30_ ( .D(n8742), .CLK(clk), .Q(arr[440]) );
  DFFPOSX1 arr_reg_10__29_ ( .D(n8741), .CLK(clk), .Q(arr[439]) );
  DFFPOSX1 arr_reg_10__28_ ( .D(n8740), .CLK(clk), .Q(arr[438]) );
  DFFPOSX1 arr_reg_10__27_ ( .D(n8739), .CLK(clk), .Q(arr[437]) );
  DFFPOSX1 arr_reg_10__26_ ( .D(n8738), .CLK(clk), .Q(arr[436]) );
  DFFPOSX1 arr_reg_10__25_ ( .D(n8737), .CLK(clk), .Q(arr[435]) );
  DFFPOSX1 arr_reg_10__24_ ( .D(n8736), .CLK(clk), .Q(arr[434]) );
  DFFPOSX1 arr_reg_10__23_ ( .D(n8735), .CLK(clk), .Q(arr[433]) );
  DFFPOSX1 arr_reg_10__22_ ( .D(n8734), .CLK(clk), .Q(arr[432]) );
  DFFPOSX1 arr_reg_10__21_ ( .D(n8733), .CLK(clk), .Q(arr[431]) );
  DFFPOSX1 arr_reg_10__20_ ( .D(n8732), .CLK(clk), .Q(arr[430]) );
  DFFPOSX1 arr_reg_10__19_ ( .D(n8731), .CLK(clk), .Q(arr[429]) );
  DFFPOSX1 arr_reg_10__18_ ( .D(n8730), .CLK(clk), .Q(arr[428]) );
  DFFPOSX1 arr_reg_10__17_ ( .D(n8729), .CLK(clk), .Q(arr[427]) );
  DFFPOSX1 arr_reg_10__16_ ( .D(n8728), .CLK(clk), .Q(arr[426]) );
  DFFPOSX1 arr_reg_10__15_ ( .D(n8727), .CLK(clk), .Q(arr[425]) );
  DFFPOSX1 arr_reg_10__14_ ( .D(n8726), .CLK(clk), .Q(arr[424]) );
  DFFPOSX1 arr_reg_10__13_ ( .D(n8725), .CLK(clk), .Q(arr[423]) );
  DFFPOSX1 arr_reg_10__12_ ( .D(n8724), .CLK(clk), .Q(arr[422]) );
  DFFPOSX1 arr_reg_10__11_ ( .D(n8723), .CLK(clk), .Q(arr[421]) );
  DFFPOSX1 arr_reg_10__10_ ( .D(n8722), .CLK(clk), .Q(arr[420]) );
  DFFPOSX1 arr_reg_10__9_ ( .D(n8721), .CLK(clk), .Q(arr[419]) );
  DFFPOSX1 arr_reg_10__8_ ( .D(n8720), .CLK(clk), .Q(arr[418]) );
  DFFPOSX1 arr_reg_10__7_ ( .D(n8719), .CLK(clk), .Q(arr[417]) );
  DFFPOSX1 arr_reg_10__6_ ( .D(n8718), .CLK(clk), .Q(arr[416]) );
  DFFPOSX1 arr_reg_10__5_ ( .D(n8717), .CLK(clk), .Q(arr[415]) );
  DFFPOSX1 arr_reg_10__4_ ( .D(n8716), .CLK(clk), .Q(arr[414]) );
  DFFPOSX1 arr_reg_10__3_ ( .D(n8715), .CLK(clk), .Q(arr[413]) );
  DFFPOSX1 arr_reg_10__2_ ( .D(n8714), .CLK(clk), .Q(arr[412]) );
  DFFPOSX1 arr_reg_10__1_ ( .D(n8713), .CLK(clk), .Q(arr[411]) );
  DFFPOSX1 arr_reg_10__0_ ( .D(n8712), .CLK(clk), .Q(arr[410]) );
  DFFPOSX1 arr_reg_9__40_ ( .D(n8711), .CLK(clk), .Q(arr[409]) );
  DFFPOSX1 arr_reg_9__39_ ( .D(n8710), .CLK(clk), .Q(arr[408]) );
  DFFPOSX1 arr_reg_9__38_ ( .D(n8709), .CLK(clk), .Q(arr[407]) );
  DFFPOSX1 arr_reg_9__37_ ( .D(n8708), .CLK(clk), .Q(arr[406]) );
  DFFPOSX1 arr_reg_9__36_ ( .D(n8707), .CLK(clk), .Q(arr[405]) );
  DFFPOSX1 arr_reg_9__35_ ( .D(n8706), .CLK(clk), .Q(arr[404]) );
  DFFPOSX1 arr_reg_9__34_ ( .D(n8705), .CLK(clk), .Q(arr[403]) );
  DFFPOSX1 arr_reg_9__33_ ( .D(n8704), .CLK(clk), .Q(arr[402]) );
  DFFPOSX1 arr_reg_9__32_ ( .D(n8703), .CLK(clk), .Q(arr[401]) );
  DFFPOSX1 arr_reg_9__31_ ( .D(n8702), .CLK(clk), .Q(arr[400]) );
  DFFPOSX1 arr_reg_9__30_ ( .D(n8701), .CLK(clk), .Q(arr[399]) );
  DFFPOSX1 arr_reg_9__29_ ( .D(n8700), .CLK(clk), .Q(arr[398]) );
  DFFPOSX1 arr_reg_9__28_ ( .D(n8699), .CLK(clk), .Q(arr[397]) );
  DFFPOSX1 arr_reg_9__27_ ( .D(n8698), .CLK(clk), .Q(arr[396]) );
  DFFPOSX1 arr_reg_9__26_ ( .D(n8697), .CLK(clk), .Q(arr[395]) );
  DFFPOSX1 arr_reg_9__25_ ( .D(n8696), .CLK(clk), .Q(arr[394]) );
  DFFPOSX1 arr_reg_9__24_ ( .D(n8695), .CLK(clk), .Q(arr[393]) );
  DFFPOSX1 arr_reg_9__23_ ( .D(n8694), .CLK(clk), .Q(arr[392]) );
  DFFPOSX1 arr_reg_9__22_ ( .D(n8693), .CLK(clk), .Q(arr[391]) );
  DFFPOSX1 arr_reg_9__21_ ( .D(n8692), .CLK(clk), .Q(arr[390]) );
  DFFPOSX1 arr_reg_9__20_ ( .D(n8691), .CLK(clk), .Q(arr[389]) );
  DFFPOSX1 arr_reg_9__19_ ( .D(n8690), .CLK(clk), .Q(arr[388]) );
  DFFPOSX1 arr_reg_9__18_ ( .D(n8689), .CLK(clk), .Q(arr[387]) );
  DFFPOSX1 arr_reg_9__17_ ( .D(n8688), .CLK(clk), .Q(arr[386]) );
  DFFPOSX1 arr_reg_9__16_ ( .D(n8687), .CLK(clk), .Q(arr[385]) );
  DFFPOSX1 arr_reg_9__15_ ( .D(n8686), .CLK(clk), .Q(arr[384]) );
  DFFPOSX1 arr_reg_9__14_ ( .D(n8685), .CLK(clk), .Q(arr[383]) );
  DFFPOSX1 arr_reg_9__13_ ( .D(n8684), .CLK(clk), .Q(arr[382]) );
  DFFPOSX1 arr_reg_9__12_ ( .D(n8683), .CLK(clk), .Q(arr[381]) );
  DFFPOSX1 arr_reg_9__11_ ( .D(n8682), .CLK(clk), .Q(arr[380]) );
  DFFPOSX1 arr_reg_9__10_ ( .D(n8681), .CLK(clk), .Q(arr[379]) );
  DFFPOSX1 arr_reg_9__9_ ( .D(n8680), .CLK(clk), .Q(arr[378]) );
  DFFPOSX1 arr_reg_9__8_ ( .D(n8679), .CLK(clk), .Q(arr[377]) );
  DFFPOSX1 arr_reg_9__7_ ( .D(n8678), .CLK(clk), .Q(arr[376]) );
  DFFPOSX1 arr_reg_9__6_ ( .D(n8677), .CLK(clk), .Q(arr[375]) );
  DFFPOSX1 arr_reg_9__5_ ( .D(n8676), .CLK(clk), .Q(arr[374]) );
  DFFPOSX1 arr_reg_9__4_ ( .D(n8675), .CLK(clk), .Q(arr[373]) );
  DFFPOSX1 arr_reg_9__3_ ( .D(n8674), .CLK(clk), .Q(arr[372]) );
  DFFPOSX1 arr_reg_9__2_ ( .D(n8673), .CLK(clk), .Q(arr[371]) );
  DFFPOSX1 arr_reg_9__1_ ( .D(n8672), .CLK(clk), .Q(arr[370]) );
  DFFPOSX1 arr_reg_9__0_ ( .D(n8671), .CLK(clk), .Q(arr[369]) );
  DFFPOSX1 arr_reg_8__40_ ( .D(n8670), .CLK(clk), .Q(arr[368]) );
  DFFPOSX1 arr_reg_8__39_ ( .D(n8669), .CLK(clk), .Q(arr[367]) );
  DFFPOSX1 arr_reg_8__38_ ( .D(n8668), .CLK(clk), .Q(arr[366]) );
  DFFPOSX1 arr_reg_8__37_ ( .D(n8667), .CLK(clk), .Q(arr[365]) );
  DFFPOSX1 arr_reg_8__36_ ( .D(n8666), .CLK(clk), .Q(arr[364]) );
  DFFPOSX1 arr_reg_8__35_ ( .D(n8665), .CLK(clk), .Q(arr[363]) );
  DFFPOSX1 arr_reg_8__34_ ( .D(n8664), .CLK(clk), .Q(arr[362]) );
  DFFPOSX1 arr_reg_8__33_ ( .D(n8663), .CLK(clk), .Q(arr[361]) );
  DFFPOSX1 arr_reg_8__32_ ( .D(n8662), .CLK(clk), .Q(arr[360]) );
  DFFPOSX1 arr_reg_8__31_ ( .D(n8661), .CLK(clk), .Q(arr[359]) );
  DFFPOSX1 arr_reg_8__30_ ( .D(n8660), .CLK(clk), .Q(arr[358]) );
  DFFPOSX1 arr_reg_8__29_ ( .D(n8659), .CLK(clk), .Q(arr[357]) );
  DFFPOSX1 arr_reg_8__28_ ( .D(n8658), .CLK(clk), .Q(arr[356]) );
  DFFPOSX1 arr_reg_8__27_ ( .D(n8657), .CLK(clk), .Q(arr[355]) );
  DFFPOSX1 arr_reg_8__26_ ( .D(n8656), .CLK(clk), .Q(arr[354]) );
  DFFPOSX1 arr_reg_8__25_ ( .D(n8655), .CLK(clk), .Q(arr[353]) );
  DFFPOSX1 arr_reg_8__24_ ( .D(n8654), .CLK(clk), .Q(arr[352]) );
  DFFPOSX1 arr_reg_8__23_ ( .D(n8653), .CLK(clk), .Q(arr[351]) );
  DFFPOSX1 arr_reg_8__22_ ( .D(n8652), .CLK(clk), .Q(arr[350]) );
  DFFPOSX1 arr_reg_8__21_ ( .D(n8651), .CLK(clk), .Q(arr[349]) );
  DFFPOSX1 arr_reg_8__20_ ( .D(n8650), .CLK(clk), .Q(arr[348]) );
  DFFPOSX1 arr_reg_8__19_ ( .D(n8649), .CLK(clk), .Q(arr[347]) );
  DFFPOSX1 arr_reg_8__18_ ( .D(n8648), .CLK(clk), .Q(arr[346]) );
  DFFPOSX1 arr_reg_8__17_ ( .D(n8647), .CLK(clk), .Q(arr[345]) );
  DFFPOSX1 arr_reg_8__16_ ( .D(n8646), .CLK(clk), .Q(arr[344]) );
  DFFPOSX1 arr_reg_8__15_ ( .D(n8645), .CLK(clk), .Q(arr[343]) );
  DFFPOSX1 arr_reg_8__14_ ( .D(n8644), .CLK(clk), .Q(arr[342]) );
  DFFPOSX1 arr_reg_8__13_ ( .D(n8643), .CLK(clk), .Q(arr[341]) );
  DFFPOSX1 arr_reg_8__12_ ( .D(n8642), .CLK(clk), .Q(arr[340]) );
  DFFPOSX1 arr_reg_8__11_ ( .D(n8641), .CLK(clk), .Q(arr[339]) );
  DFFPOSX1 arr_reg_8__10_ ( .D(n8640), .CLK(clk), .Q(arr[338]) );
  DFFPOSX1 arr_reg_8__9_ ( .D(n8639), .CLK(clk), .Q(arr[337]) );
  DFFPOSX1 arr_reg_8__8_ ( .D(n8638), .CLK(clk), .Q(arr[336]) );
  DFFPOSX1 arr_reg_8__7_ ( .D(n8637), .CLK(clk), .Q(arr[335]) );
  DFFPOSX1 arr_reg_8__6_ ( .D(n8636), .CLK(clk), .Q(arr[334]) );
  DFFPOSX1 arr_reg_8__5_ ( .D(n8635), .CLK(clk), .Q(arr[333]) );
  DFFPOSX1 arr_reg_8__4_ ( .D(n8634), .CLK(clk), .Q(arr[332]) );
  DFFPOSX1 arr_reg_8__3_ ( .D(n8633), .CLK(clk), .Q(arr[331]) );
  DFFPOSX1 arr_reg_8__2_ ( .D(n8632), .CLK(clk), .Q(arr[330]) );
  DFFPOSX1 arr_reg_8__1_ ( .D(n8631), .CLK(clk), .Q(arr[329]) );
  DFFPOSX1 arr_reg_8__0_ ( .D(n8630), .CLK(clk), .Q(arr[328]) );
  DFFPOSX1 arr_reg_7__40_ ( .D(n8629), .CLK(clk), .Q(arr[327]) );
  DFFPOSX1 arr_reg_7__39_ ( .D(n8628), .CLK(clk), .Q(arr[326]) );
  DFFPOSX1 arr_reg_7__38_ ( .D(n8627), .CLK(clk), .Q(arr[325]) );
  DFFPOSX1 arr_reg_7__37_ ( .D(n8626), .CLK(clk), .Q(arr[324]) );
  DFFPOSX1 arr_reg_7__36_ ( .D(n8625), .CLK(clk), .Q(arr[323]) );
  DFFPOSX1 arr_reg_7__35_ ( .D(n8624), .CLK(clk), .Q(arr[322]) );
  DFFPOSX1 arr_reg_7__34_ ( .D(n8623), .CLK(clk), .Q(arr[321]) );
  DFFPOSX1 arr_reg_7__33_ ( .D(n8622), .CLK(clk), .Q(arr[320]) );
  DFFPOSX1 arr_reg_7__32_ ( .D(n8621), .CLK(clk), .Q(arr[319]) );
  DFFPOSX1 arr_reg_7__31_ ( .D(n8620), .CLK(clk), .Q(arr[318]) );
  DFFPOSX1 arr_reg_7__30_ ( .D(n8619), .CLK(clk), .Q(arr[317]) );
  DFFPOSX1 arr_reg_7__29_ ( .D(n8618), .CLK(clk), .Q(arr[316]) );
  DFFPOSX1 arr_reg_7__28_ ( .D(n8617), .CLK(clk), .Q(arr[315]) );
  DFFPOSX1 arr_reg_7__27_ ( .D(n8616), .CLK(clk), .Q(arr[314]) );
  DFFPOSX1 arr_reg_7__26_ ( .D(n8615), .CLK(clk), .Q(arr[313]) );
  DFFPOSX1 arr_reg_7__25_ ( .D(n8614), .CLK(clk), .Q(arr[312]) );
  DFFPOSX1 arr_reg_7__24_ ( .D(n8613), .CLK(clk), .Q(arr[311]) );
  DFFPOSX1 arr_reg_7__23_ ( .D(n8612), .CLK(clk), .Q(arr[310]) );
  DFFPOSX1 arr_reg_7__22_ ( .D(n8611), .CLK(clk), .Q(arr[309]) );
  DFFPOSX1 arr_reg_7__21_ ( .D(n8610), .CLK(clk), .Q(arr[308]) );
  DFFPOSX1 arr_reg_7__20_ ( .D(n8609), .CLK(clk), .Q(arr[307]) );
  DFFPOSX1 arr_reg_7__19_ ( .D(n8608), .CLK(clk), .Q(arr[306]) );
  DFFPOSX1 arr_reg_7__18_ ( .D(n8607), .CLK(clk), .Q(arr[305]) );
  DFFPOSX1 arr_reg_7__17_ ( .D(n8606), .CLK(clk), .Q(arr[304]) );
  DFFPOSX1 arr_reg_7__16_ ( .D(n8605), .CLK(clk), .Q(arr[303]) );
  DFFPOSX1 arr_reg_7__15_ ( .D(n8604), .CLK(clk), .Q(arr[302]) );
  DFFPOSX1 arr_reg_7__14_ ( .D(n8603), .CLK(clk), .Q(arr[301]) );
  DFFPOSX1 arr_reg_7__13_ ( .D(n8602), .CLK(clk), .Q(arr[300]) );
  DFFPOSX1 arr_reg_7__12_ ( .D(n8601), .CLK(clk), .Q(arr[299]) );
  DFFPOSX1 arr_reg_7__11_ ( .D(n8600), .CLK(clk), .Q(arr[298]) );
  DFFPOSX1 arr_reg_7__10_ ( .D(n8599), .CLK(clk), .Q(arr[297]) );
  DFFPOSX1 arr_reg_7__9_ ( .D(n8598), .CLK(clk), .Q(arr[296]) );
  DFFPOSX1 arr_reg_7__8_ ( .D(n8597), .CLK(clk), .Q(arr[295]) );
  DFFPOSX1 arr_reg_7__7_ ( .D(n8596), .CLK(clk), .Q(arr[294]) );
  DFFPOSX1 arr_reg_7__6_ ( .D(n8595), .CLK(clk), .Q(arr[293]) );
  DFFPOSX1 arr_reg_7__5_ ( .D(n8594), .CLK(clk), .Q(arr[292]) );
  DFFPOSX1 arr_reg_7__4_ ( .D(n8593), .CLK(clk), .Q(arr[291]) );
  DFFPOSX1 arr_reg_7__3_ ( .D(n8592), .CLK(clk), .Q(arr[290]) );
  DFFPOSX1 arr_reg_7__2_ ( .D(n8591), .CLK(clk), .Q(arr[289]) );
  DFFPOSX1 arr_reg_7__1_ ( .D(n8590), .CLK(clk), .Q(arr[288]) );
  DFFPOSX1 arr_reg_7__0_ ( .D(n8589), .CLK(clk), .Q(arr[287]) );
  DFFPOSX1 arr_reg_6__40_ ( .D(n8588), .CLK(clk), .Q(arr[286]) );
  DFFPOSX1 arr_reg_6__39_ ( .D(n8587), .CLK(clk), .Q(arr[285]) );
  DFFPOSX1 arr_reg_6__38_ ( .D(n8586), .CLK(clk), .Q(arr[284]) );
  DFFPOSX1 arr_reg_6__37_ ( .D(n8585), .CLK(clk), .Q(arr[283]) );
  DFFPOSX1 arr_reg_6__36_ ( .D(n8584), .CLK(clk), .Q(arr[282]) );
  DFFPOSX1 arr_reg_6__35_ ( .D(n8583), .CLK(clk), .Q(arr[281]) );
  DFFPOSX1 arr_reg_6__34_ ( .D(n8582), .CLK(clk), .Q(arr[280]) );
  DFFPOSX1 arr_reg_6__33_ ( .D(n8581), .CLK(clk), .Q(arr[279]) );
  DFFPOSX1 arr_reg_6__32_ ( .D(n8580), .CLK(clk), .Q(arr[278]) );
  DFFPOSX1 arr_reg_6__31_ ( .D(n8579), .CLK(clk), .Q(arr[277]) );
  DFFPOSX1 arr_reg_6__30_ ( .D(n8578), .CLK(clk), .Q(arr[276]) );
  DFFPOSX1 arr_reg_6__29_ ( .D(n8577), .CLK(clk), .Q(arr[275]) );
  DFFPOSX1 arr_reg_6__28_ ( .D(n8576), .CLK(clk), .Q(arr[274]) );
  DFFPOSX1 arr_reg_6__27_ ( .D(n8575), .CLK(clk), .Q(arr[273]) );
  DFFPOSX1 arr_reg_6__26_ ( .D(n8574), .CLK(clk), .Q(arr[272]) );
  DFFPOSX1 arr_reg_6__25_ ( .D(n8573), .CLK(clk), .Q(arr[271]) );
  DFFPOSX1 arr_reg_6__24_ ( .D(n8572), .CLK(clk), .Q(arr[270]) );
  DFFPOSX1 arr_reg_6__23_ ( .D(n8571), .CLK(clk), .Q(arr[269]) );
  DFFPOSX1 arr_reg_6__22_ ( .D(n8570), .CLK(clk), .Q(arr[268]) );
  DFFPOSX1 arr_reg_6__21_ ( .D(n8569), .CLK(clk), .Q(arr[267]) );
  DFFPOSX1 arr_reg_6__20_ ( .D(n8568), .CLK(clk), .Q(arr[266]) );
  DFFPOSX1 arr_reg_6__19_ ( .D(n8567), .CLK(clk), .Q(arr[265]) );
  DFFPOSX1 arr_reg_6__18_ ( .D(n8566), .CLK(clk), .Q(arr[264]) );
  DFFPOSX1 arr_reg_6__17_ ( .D(n8565), .CLK(clk), .Q(arr[263]) );
  DFFPOSX1 arr_reg_6__16_ ( .D(n8564), .CLK(clk), .Q(arr[262]) );
  DFFPOSX1 arr_reg_6__15_ ( .D(n8563), .CLK(clk), .Q(arr[261]) );
  DFFPOSX1 arr_reg_6__14_ ( .D(n8562), .CLK(clk), .Q(arr[260]) );
  DFFPOSX1 arr_reg_6__13_ ( .D(n8561), .CLK(clk), .Q(arr[259]) );
  DFFPOSX1 arr_reg_6__12_ ( .D(n8560), .CLK(clk), .Q(arr[258]) );
  DFFPOSX1 arr_reg_6__11_ ( .D(n8559), .CLK(clk), .Q(arr[257]) );
  DFFPOSX1 arr_reg_6__10_ ( .D(n8558), .CLK(clk), .Q(arr[256]) );
  DFFPOSX1 arr_reg_6__9_ ( .D(n8557), .CLK(clk), .Q(arr[255]) );
  DFFPOSX1 arr_reg_6__8_ ( .D(n8556), .CLK(clk), .Q(arr[254]) );
  DFFPOSX1 arr_reg_6__7_ ( .D(n8555), .CLK(clk), .Q(arr[253]) );
  DFFPOSX1 arr_reg_6__6_ ( .D(n8554), .CLK(clk), .Q(arr[252]) );
  DFFPOSX1 arr_reg_6__5_ ( .D(n8553), .CLK(clk), .Q(arr[251]) );
  DFFPOSX1 arr_reg_6__4_ ( .D(n8552), .CLK(clk), .Q(arr[250]) );
  DFFPOSX1 arr_reg_6__3_ ( .D(n8551), .CLK(clk), .Q(arr[249]) );
  DFFPOSX1 arr_reg_6__2_ ( .D(n8550), .CLK(clk), .Q(arr[248]) );
  DFFPOSX1 arr_reg_6__1_ ( .D(n8549), .CLK(clk), .Q(arr[247]) );
  DFFPOSX1 arr_reg_6__0_ ( .D(n8548), .CLK(clk), .Q(arr[246]) );
  DFFPOSX1 arr_reg_5__40_ ( .D(n8547), .CLK(clk), .Q(arr[245]) );
  DFFPOSX1 arr_reg_5__39_ ( .D(n8546), .CLK(clk), .Q(arr[244]) );
  DFFPOSX1 arr_reg_5__38_ ( .D(n8545), .CLK(clk), .Q(arr[243]) );
  DFFPOSX1 arr_reg_5__37_ ( .D(n8544), .CLK(clk), .Q(arr[242]) );
  DFFPOSX1 arr_reg_5__36_ ( .D(n8543), .CLK(clk), .Q(arr[241]) );
  DFFPOSX1 arr_reg_5__35_ ( .D(n8542), .CLK(clk), .Q(arr[240]) );
  DFFPOSX1 arr_reg_5__34_ ( .D(n8541), .CLK(clk), .Q(arr[239]) );
  DFFPOSX1 arr_reg_5__33_ ( .D(n8540), .CLK(clk), .Q(arr[238]) );
  DFFPOSX1 arr_reg_5__32_ ( .D(n8539), .CLK(clk), .Q(arr[237]) );
  DFFPOSX1 arr_reg_5__31_ ( .D(n8538), .CLK(clk), .Q(arr[236]) );
  DFFPOSX1 arr_reg_5__30_ ( .D(n8537), .CLK(clk), .Q(arr[235]) );
  DFFPOSX1 arr_reg_5__29_ ( .D(n8536), .CLK(clk), .Q(arr[234]) );
  DFFPOSX1 arr_reg_5__28_ ( .D(n8535), .CLK(clk), .Q(arr[233]) );
  DFFPOSX1 arr_reg_5__27_ ( .D(n8534), .CLK(clk), .Q(arr[232]) );
  DFFPOSX1 arr_reg_5__26_ ( .D(n8533), .CLK(clk), .Q(arr[231]) );
  DFFPOSX1 arr_reg_5__25_ ( .D(n8532), .CLK(clk), .Q(arr[230]) );
  DFFPOSX1 arr_reg_5__24_ ( .D(n8531), .CLK(clk), .Q(arr[229]) );
  DFFPOSX1 arr_reg_5__23_ ( .D(n8530), .CLK(clk), .Q(arr[228]) );
  DFFPOSX1 arr_reg_5__22_ ( .D(n8529), .CLK(clk), .Q(arr[227]) );
  DFFPOSX1 arr_reg_5__21_ ( .D(n8528), .CLK(clk), .Q(arr[226]) );
  DFFPOSX1 arr_reg_5__20_ ( .D(n8527), .CLK(clk), .Q(arr[225]) );
  DFFPOSX1 arr_reg_5__19_ ( .D(n8526), .CLK(clk), .Q(arr[224]) );
  DFFPOSX1 arr_reg_5__18_ ( .D(n8525), .CLK(clk), .Q(arr[223]) );
  DFFPOSX1 arr_reg_5__17_ ( .D(n8524), .CLK(clk), .Q(arr[222]) );
  DFFPOSX1 arr_reg_5__16_ ( .D(n8523), .CLK(clk), .Q(arr[221]) );
  DFFPOSX1 arr_reg_5__15_ ( .D(n8522), .CLK(clk), .Q(arr[220]) );
  DFFPOSX1 arr_reg_5__14_ ( .D(n8521), .CLK(clk), .Q(arr[219]) );
  DFFPOSX1 arr_reg_5__13_ ( .D(n8520), .CLK(clk), .Q(arr[218]) );
  DFFPOSX1 arr_reg_5__12_ ( .D(n8519), .CLK(clk), .Q(arr[217]) );
  DFFPOSX1 arr_reg_5__11_ ( .D(n8518), .CLK(clk), .Q(arr[216]) );
  DFFPOSX1 arr_reg_5__10_ ( .D(n8517), .CLK(clk), .Q(arr[215]) );
  DFFPOSX1 arr_reg_5__9_ ( .D(n8516), .CLK(clk), .Q(arr[214]) );
  DFFPOSX1 arr_reg_5__8_ ( .D(n8515), .CLK(clk), .Q(arr[213]) );
  DFFPOSX1 arr_reg_5__7_ ( .D(n8514), .CLK(clk), .Q(arr[212]) );
  DFFPOSX1 arr_reg_5__6_ ( .D(n8513), .CLK(clk), .Q(arr[211]) );
  DFFPOSX1 arr_reg_5__5_ ( .D(n8512), .CLK(clk), .Q(arr[210]) );
  DFFPOSX1 arr_reg_5__4_ ( .D(n8511), .CLK(clk), .Q(arr[209]) );
  DFFPOSX1 arr_reg_5__3_ ( .D(n8510), .CLK(clk), .Q(arr[208]) );
  DFFPOSX1 arr_reg_5__2_ ( .D(n8509), .CLK(clk), .Q(arr[207]) );
  DFFPOSX1 arr_reg_5__1_ ( .D(n8508), .CLK(clk), .Q(arr[206]) );
  DFFPOSX1 arr_reg_5__0_ ( .D(n8507), .CLK(clk), .Q(arr[205]) );
  DFFPOSX1 arr_reg_4__40_ ( .D(n8506), .CLK(clk), .Q(arr[204]) );
  DFFPOSX1 arr_reg_4__39_ ( .D(n8505), .CLK(clk), .Q(arr[203]) );
  DFFPOSX1 arr_reg_4__38_ ( .D(n8504), .CLK(clk), .Q(arr[202]) );
  DFFPOSX1 arr_reg_4__37_ ( .D(n8503), .CLK(clk), .Q(arr[201]) );
  DFFPOSX1 arr_reg_4__36_ ( .D(n8502), .CLK(clk), .Q(arr[200]) );
  DFFPOSX1 arr_reg_4__35_ ( .D(n8501), .CLK(clk), .Q(arr[199]) );
  DFFPOSX1 arr_reg_4__34_ ( .D(n8500), .CLK(clk), .Q(arr[198]) );
  DFFPOSX1 arr_reg_4__33_ ( .D(n8499), .CLK(clk), .Q(arr[197]) );
  DFFPOSX1 arr_reg_4__32_ ( .D(n8498), .CLK(clk), .Q(arr[196]) );
  DFFPOSX1 arr_reg_4__31_ ( .D(n8497), .CLK(clk), .Q(arr[195]) );
  DFFPOSX1 arr_reg_4__30_ ( .D(n8496), .CLK(clk), .Q(arr[194]) );
  DFFPOSX1 arr_reg_4__29_ ( .D(n8495), .CLK(clk), .Q(arr[193]) );
  DFFPOSX1 arr_reg_4__28_ ( .D(n8494), .CLK(clk), .Q(arr[192]) );
  DFFPOSX1 arr_reg_4__27_ ( .D(n8493), .CLK(clk), .Q(arr[191]) );
  DFFPOSX1 arr_reg_4__26_ ( .D(n8492), .CLK(clk), .Q(arr[190]) );
  DFFPOSX1 arr_reg_4__25_ ( .D(n8491), .CLK(clk), .Q(arr[189]) );
  DFFPOSX1 arr_reg_4__24_ ( .D(n8490), .CLK(clk), .Q(arr[188]) );
  DFFPOSX1 arr_reg_4__23_ ( .D(n8489), .CLK(clk), .Q(arr[187]) );
  DFFPOSX1 arr_reg_4__22_ ( .D(n8488), .CLK(clk), .Q(arr[186]) );
  DFFPOSX1 arr_reg_4__21_ ( .D(n8487), .CLK(clk), .Q(arr[185]) );
  DFFPOSX1 arr_reg_4__20_ ( .D(n8486), .CLK(clk), .Q(arr[184]) );
  DFFPOSX1 arr_reg_4__19_ ( .D(n8485), .CLK(clk), .Q(arr[183]) );
  DFFPOSX1 arr_reg_4__18_ ( .D(n8484), .CLK(clk), .Q(arr[182]) );
  DFFPOSX1 arr_reg_4__17_ ( .D(n8483), .CLK(clk), .Q(arr[181]) );
  DFFPOSX1 arr_reg_4__16_ ( .D(n8482), .CLK(clk), .Q(arr[180]) );
  DFFPOSX1 arr_reg_4__15_ ( .D(n8481), .CLK(clk), .Q(arr[179]) );
  DFFPOSX1 arr_reg_4__14_ ( .D(n8480), .CLK(clk), .Q(arr[178]) );
  DFFPOSX1 arr_reg_4__13_ ( .D(n8479), .CLK(clk), .Q(arr[177]) );
  DFFPOSX1 arr_reg_4__12_ ( .D(n8478), .CLK(clk), .Q(arr[176]) );
  DFFPOSX1 arr_reg_4__11_ ( .D(n8477), .CLK(clk), .Q(arr[175]) );
  DFFPOSX1 arr_reg_4__10_ ( .D(n8476), .CLK(clk), .Q(arr[174]) );
  DFFPOSX1 arr_reg_4__9_ ( .D(n8475), .CLK(clk), .Q(arr[173]) );
  DFFPOSX1 arr_reg_4__8_ ( .D(n8474), .CLK(clk), .Q(arr[172]) );
  DFFPOSX1 arr_reg_4__7_ ( .D(n8473), .CLK(clk), .Q(arr[171]) );
  DFFPOSX1 arr_reg_4__6_ ( .D(n8472), .CLK(clk), .Q(arr[170]) );
  DFFPOSX1 arr_reg_4__5_ ( .D(n8471), .CLK(clk), .Q(arr[169]) );
  DFFPOSX1 arr_reg_4__4_ ( .D(n8470), .CLK(clk), .Q(arr[168]) );
  DFFPOSX1 arr_reg_4__3_ ( .D(n8469), .CLK(clk), .Q(arr[167]) );
  DFFPOSX1 arr_reg_4__2_ ( .D(n8468), .CLK(clk), .Q(arr[166]) );
  DFFPOSX1 arr_reg_4__1_ ( .D(n8467), .CLK(clk), .Q(arr[165]) );
  DFFPOSX1 arr_reg_4__0_ ( .D(n8466), .CLK(clk), .Q(arr[164]) );
  DFFPOSX1 arr_reg_3__40_ ( .D(n8465), .CLK(clk), .Q(arr[163]) );
  DFFPOSX1 arr_reg_3__39_ ( .D(n8464), .CLK(clk), .Q(arr[162]) );
  DFFPOSX1 arr_reg_3__38_ ( .D(n8463), .CLK(clk), .Q(arr[161]) );
  DFFPOSX1 arr_reg_3__37_ ( .D(n8462), .CLK(clk), .Q(arr[160]) );
  DFFPOSX1 arr_reg_3__36_ ( .D(n8461), .CLK(clk), .Q(arr[159]) );
  DFFPOSX1 arr_reg_3__35_ ( .D(n8460), .CLK(clk), .Q(arr[158]) );
  DFFPOSX1 arr_reg_3__34_ ( .D(n8459), .CLK(clk), .Q(arr[157]) );
  DFFPOSX1 arr_reg_3__33_ ( .D(n8458), .CLK(clk), .Q(arr[156]) );
  DFFPOSX1 arr_reg_3__32_ ( .D(n8457), .CLK(clk), .Q(arr[155]) );
  DFFPOSX1 arr_reg_3__31_ ( .D(n8456), .CLK(clk), .Q(arr[154]) );
  DFFPOSX1 arr_reg_3__30_ ( .D(n8455), .CLK(clk), .Q(arr[153]) );
  DFFPOSX1 arr_reg_3__29_ ( .D(n8454), .CLK(clk), .Q(arr[152]) );
  DFFPOSX1 arr_reg_3__28_ ( .D(n8453), .CLK(clk), .Q(arr[151]) );
  DFFPOSX1 arr_reg_3__27_ ( .D(n8452), .CLK(clk), .Q(arr[150]) );
  DFFPOSX1 arr_reg_3__26_ ( .D(n8451), .CLK(clk), .Q(arr[149]) );
  DFFPOSX1 arr_reg_3__25_ ( .D(n8450), .CLK(clk), .Q(arr[148]) );
  DFFPOSX1 arr_reg_3__24_ ( .D(n8449), .CLK(clk), .Q(arr[147]) );
  DFFPOSX1 arr_reg_3__23_ ( .D(n8448), .CLK(clk), .Q(arr[146]) );
  DFFPOSX1 arr_reg_3__22_ ( .D(n8447), .CLK(clk), .Q(arr[145]) );
  DFFPOSX1 arr_reg_3__21_ ( .D(n8446), .CLK(clk), .Q(arr[144]) );
  DFFPOSX1 arr_reg_3__20_ ( .D(n8445), .CLK(clk), .Q(arr[143]) );
  DFFPOSX1 arr_reg_3__19_ ( .D(n8444), .CLK(clk), .Q(arr[142]) );
  DFFPOSX1 arr_reg_3__18_ ( .D(n8443), .CLK(clk), .Q(arr[141]) );
  DFFPOSX1 arr_reg_3__17_ ( .D(n8442), .CLK(clk), .Q(arr[140]) );
  DFFPOSX1 arr_reg_3__16_ ( .D(n8441), .CLK(clk), .Q(arr[139]) );
  DFFPOSX1 arr_reg_3__15_ ( .D(n8440), .CLK(clk), .Q(arr[138]) );
  DFFPOSX1 arr_reg_3__14_ ( .D(n8439), .CLK(clk), .Q(arr[137]) );
  DFFPOSX1 arr_reg_3__13_ ( .D(n8438), .CLK(clk), .Q(arr[136]) );
  DFFPOSX1 arr_reg_3__12_ ( .D(n8437), .CLK(clk), .Q(arr[135]) );
  DFFPOSX1 arr_reg_3__11_ ( .D(n8436), .CLK(clk), .Q(arr[134]) );
  DFFPOSX1 arr_reg_3__10_ ( .D(n8435), .CLK(clk), .Q(arr[133]) );
  DFFPOSX1 arr_reg_3__9_ ( .D(n8434), .CLK(clk), .Q(arr[132]) );
  DFFPOSX1 arr_reg_3__8_ ( .D(n8433), .CLK(clk), .Q(arr[131]) );
  DFFPOSX1 arr_reg_3__7_ ( .D(n8432), .CLK(clk), .Q(arr[130]) );
  DFFPOSX1 arr_reg_3__6_ ( .D(n8431), .CLK(clk), .Q(arr[129]) );
  DFFPOSX1 arr_reg_3__5_ ( .D(n8430), .CLK(clk), .Q(arr[128]) );
  DFFPOSX1 arr_reg_3__4_ ( .D(n8429), .CLK(clk), .Q(arr[127]) );
  DFFPOSX1 arr_reg_3__3_ ( .D(n8428), .CLK(clk), .Q(arr[126]) );
  DFFPOSX1 arr_reg_3__2_ ( .D(n8427), .CLK(clk), .Q(arr[125]) );
  DFFPOSX1 arr_reg_3__1_ ( .D(n8426), .CLK(clk), .Q(arr[124]) );
  DFFPOSX1 arr_reg_3__0_ ( .D(n8425), .CLK(clk), .Q(arr[123]) );
  DFFPOSX1 arr_reg_2__40_ ( .D(n8424), .CLK(clk), .Q(arr[122]) );
  DFFPOSX1 arr_reg_2__39_ ( .D(n8423), .CLK(clk), .Q(arr[121]) );
  DFFPOSX1 arr_reg_2__38_ ( .D(n8422), .CLK(clk), .Q(arr[120]) );
  DFFPOSX1 arr_reg_2__37_ ( .D(n8421), .CLK(clk), .Q(arr[119]) );
  DFFPOSX1 arr_reg_2__36_ ( .D(n8420), .CLK(clk), .Q(arr[118]) );
  DFFPOSX1 arr_reg_2__35_ ( .D(n8419), .CLK(clk), .Q(arr[117]) );
  DFFPOSX1 arr_reg_2__34_ ( .D(n8418), .CLK(clk), .Q(arr[116]) );
  DFFPOSX1 arr_reg_2__33_ ( .D(n8417), .CLK(clk), .Q(arr[115]) );
  DFFPOSX1 arr_reg_2__32_ ( .D(n8416), .CLK(clk), .Q(arr[114]) );
  DFFPOSX1 arr_reg_2__31_ ( .D(n8415), .CLK(clk), .Q(arr[113]) );
  DFFPOSX1 arr_reg_2__30_ ( .D(n8414), .CLK(clk), .Q(arr[112]) );
  DFFPOSX1 arr_reg_2__29_ ( .D(n8413), .CLK(clk), .Q(arr[111]) );
  DFFPOSX1 arr_reg_2__28_ ( .D(n8412), .CLK(clk), .Q(arr[110]) );
  DFFPOSX1 arr_reg_2__27_ ( .D(n8411), .CLK(clk), .Q(arr[109]) );
  DFFPOSX1 arr_reg_2__26_ ( .D(n8410), .CLK(clk), .Q(arr[108]) );
  DFFPOSX1 arr_reg_2__25_ ( .D(n8409), .CLK(clk), .Q(arr[107]) );
  DFFPOSX1 arr_reg_2__24_ ( .D(n8408), .CLK(clk), .Q(arr[106]) );
  DFFPOSX1 arr_reg_2__23_ ( .D(n8407), .CLK(clk), .Q(arr[105]) );
  DFFPOSX1 arr_reg_2__22_ ( .D(n8406), .CLK(clk), .Q(arr[104]) );
  DFFPOSX1 arr_reg_2__21_ ( .D(n8405), .CLK(clk), .Q(arr[103]) );
  DFFPOSX1 arr_reg_2__20_ ( .D(n8404), .CLK(clk), .Q(arr[102]) );
  DFFPOSX1 arr_reg_2__19_ ( .D(n8403), .CLK(clk), .Q(arr[101]) );
  DFFPOSX1 arr_reg_2__18_ ( .D(n8402), .CLK(clk), .Q(arr[100]) );
  DFFPOSX1 arr_reg_2__17_ ( .D(n8401), .CLK(clk), .Q(arr[99]) );
  DFFPOSX1 arr_reg_2__16_ ( .D(n8400), .CLK(clk), .Q(arr[98]) );
  DFFPOSX1 arr_reg_2__15_ ( .D(n8399), .CLK(clk), .Q(arr[97]) );
  DFFPOSX1 arr_reg_2__14_ ( .D(n8398), .CLK(clk), .Q(arr[96]) );
  DFFPOSX1 arr_reg_2__13_ ( .D(n8397), .CLK(clk), .Q(arr[95]) );
  DFFPOSX1 arr_reg_2__12_ ( .D(n8396), .CLK(clk), .Q(arr[94]) );
  DFFPOSX1 arr_reg_2__11_ ( .D(n8395), .CLK(clk), .Q(arr[93]) );
  DFFPOSX1 arr_reg_2__10_ ( .D(n8394), .CLK(clk), .Q(arr[92]) );
  DFFPOSX1 arr_reg_2__9_ ( .D(n8393), .CLK(clk), .Q(arr[91]) );
  DFFPOSX1 arr_reg_2__8_ ( .D(n8392), .CLK(clk), .Q(arr[90]) );
  DFFPOSX1 arr_reg_2__7_ ( .D(n8391), .CLK(clk), .Q(arr[89]) );
  DFFPOSX1 arr_reg_2__6_ ( .D(n8390), .CLK(clk), .Q(arr[88]) );
  DFFPOSX1 arr_reg_2__5_ ( .D(n8389), .CLK(clk), .Q(arr[87]) );
  DFFPOSX1 arr_reg_2__4_ ( .D(n8388), .CLK(clk), .Q(arr[86]) );
  DFFPOSX1 arr_reg_2__3_ ( .D(n8387), .CLK(clk), .Q(arr[85]) );
  DFFPOSX1 arr_reg_2__2_ ( .D(n8386), .CLK(clk), .Q(arr[84]) );
  DFFPOSX1 arr_reg_2__1_ ( .D(n8385), .CLK(clk), .Q(arr[83]) );
  DFFPOSX1 arr_reg_2__0_ ( .D(n8384), .CLK(clk), .Q(arr[82]) );
  DFFPOSX1 arr_reg_1__40_ ( .D(n8383), .CLK(clk), .Q(arr[81]) );
  DFFPOSX1 arr_reg_1__39_ ( .D(n8382), .CLK(clk), .Q(arr[80]) );
  DFFPOSX1 arr_reg_1__38_ ( .D(n8381), .CLK(clk), .Q(arr[79]) );
  DFFPOSX1 arr_reg_1__37_ ( .D(n8380), .CLK(clk), .Q(arr[78]) );
  DFFPOSX1 arr_reg_1__36_ ( .D(n8379), .CLK(clk), .Q(arr[77]) );
  DFFPOSX1 arr_reg_1__35_ ( .D(n8378), .CLK(clk), .Q(arr[76]) );
  DFFPOSX1 arr_reg_1__34_ ( .D(n8377), .CLK(clk), .Q(arr[75]) );
  DFFPOSX1 arr_reg_1__33_ ( .D(n8376), .CLK(clk), .Q(arr[74]) );
  DFFPOSX1 arr_reg_1__32_ ( .D(n8375), .CLK(clk), .Q(arr[73]) );
  DFFPOSX1 arr_reg_1__31_ ( .D(n8374), .CLK(clk), .Q(arr[72]) );
  DFFPOSX1 arr_reg_1__30_ ( .D(n8373), .CLK(clk), .Q(arr[71]) );
  DFFPOSX1 arr_reg_1__29_ ( .D(n8372), .CLK(clk), .Q(arr[70]) );
  DFFPOSX1 arr_reg_1__28_ ( .D(n8371), .CLK(clk), .Q(arr[69]) );
  DFFPOSX1 arr_reg_1__27_ ( .D(n8370), .CLK(clk), .Q(arr[68]) );
  DFFPOSX1 arr_reg_1__26_ ( .D(n8369), .CLK(clk), .Q(arr[67]) );
  DFFPOSX1 arr_reg_1__25_ ( .D(n8368), .CLK(clk), .Q(arr[66]) );
  DFFPOSX1 arr_reg_1__24_ ( .D(n8367), .CLK(clk), .Q(arr[65]) );
  DFFPOSX1 arr_reg_1__23_ ( .D(n8366), .CLK(clk), .Q(arr[64]) );
  DFFPOSX1 arr_reg_1__22_ ( .D(n8365), .CLK(clk), .Q(arr[63]) );
  DFFPOSX1 arr_reg_1__21_ ( .D(n8364), .CLK(clk), .Q(arr[62]) );
  DFFPOSX1 arr_reg_1__20_ ( .D(n8363), .CLK(clk), .Q(arr[61]) );
  DFFPOSX1 arr_reg_1__19_ ( .D(n8362), .CLK(clk), .Q(arr[60]) );
  DFFPOSX1 arr_reg_1__18_ ( .D(n8361), .CLK(clk), .Q(arr[59]) );
  DFFPOSX1 arr_reg_1__17_ ( .D(n8360), .CLK(clk), .Q(arr[58]) );
  DFFPOSX1 arr_reg_1__16_ ( .D(n8359), .CLK(clk), .Q(arr[57]) );
  DFFPOSX1 arr_reg_1__15_ ( .D(n8358), .CLK(clk), .Q(arr[56]) );
  DFFPOSX1 arr_reg_1__14_ ( .D(n8357), .CLK(clk), .Q(arr[55]) );
  DFFPOSX1 arr_reg_1__13_ ( .D(n8356), .CLK(clk), .Q(arr[54]) );
  DFFPOSX1 arr_reg_1__12_ ( .D(n8355), .CLK(clk), .Q(arr[53]) );
  DFFPOSX1 arr_reg_1__11_ ( .D(n8354), .CLK(clk), .Q(arr[52]) );
  DFFPOSX1 arr_reg_1__10_ ( .D(n8353), .CLK(clk), .Q(arr[51]) );
  DFFPOSX1 arr_reg_1__9_ ( .D(n8352), .CLK(clk), .Q(arr[50]) );
  DFFPOSX1 arr_reg_1__8_ ( .D(n8351), .CLK(clk), .Q(arr[49]) );
  DFFPOSX1 arr_reg_1__7_ ( .D(n8350), .CLK(clk), .Q(arr[48]) );
  DFFPOSX1 arr_reg_1__6_ ( .D(n8349), .CLK(clk), .Q(arr[47]) );
  DFFPOSX1 arr_reg_1__5_ ( .D(n8348), .CLK(clk), .Q(arr[46]) );
  DFFPOSX1 arr_reg_1__4_ ( .D(n8347), .CLK(clk), .Q(arr[45]) );
  DFFPOSX1 arr_reg_1__3_ ( .D(n8346), .CLK(clk), .Q(arr[44]) );
  DFFPOSX1 arr_reg_1__2_ ( .D(n8345), .CLK(clk), .Q(arr[43]) );
  DFFPOSX1 arr_reg_1__1_ ( .D(n8344), .CLK(clk), .Q(arr[42]) );
  DFFPOSX1 arr_reg_1__0_ ( .D(n8343), .CLK(clk), .Q(arr[41]) );
  DFFPOSX1 arr_reg_0__40_ ( .D(n8342), .CLK(clk), .Q(arr[40]) );
  DFFPOSX1 arr_reg_0__39_ ( .D(n8341), .CLK(clk), .Q(arr[39]) );
  DFFPOSX1 arr_reg_0__38_ ( .D(n8340), .CLK(clk), .Q(arr[38]) );
  DFFPOSX1 arr_reg_0__37_ ( .D(n8339), .CLK(clk), .Q(arr[37]) );
  DFFPOSX1 arr_reg_0__36_ ( .D(n8338), .CLK(clk), .Q(arr[36]) );
  DFFPOSX1 arr_reg_0__35_ ( .D(n8337), .CLK(clk), .Q(arr[35]) );
  DFFPOSX1 arr_reg_0__34_ ( .D(n8336), .CLK(clk), .Q(arr[34]) );
  DFFPOSX1 arr_reg_0__33_ ( .D(n8335), .CLK(clk), .Q(arr[33]) );
  DFFPOSX1 arr_reg_0__32_ ( .D(n8334), .CLK(clk), .Q(arr[32]) );
  DFFPOSX1 arr_reg_0__31_ ( .D(n8333), .CLK(clk), .Q(arr[31]) );
  DFFPOSX1 arr_reg_0__30_ ( .D(n8332), .CLK(clk), .Q(arr[30]) );
  DFFPOSX1 arr_reg_0__29_ ( .D(n8331), .CLK(clk), .Q(arr[29]) );
  DFFPOSX1 arr_reg_0__28_ ( .D(n8330), .CLK(clk), .Q(arr[28]) );
  DFFPOSX1 arr_reg_0__27_ ( .D(n8329), .CLK(clk), .Q(arr[27]) );
  DFFPOSX1 arr_reg_0__26_ ( .D(n8328), .CLK(clk), .Q(arr[26]) );
  DFFPOSX1 arr_reg_0__25_ ( .D(n8327), .CLK(clk), .Q(arr[25]) );
  DFFPOSX1 arr_reg_0__24_ ( .D(n8326), .CLK(clk), .Q(arr[24]) );
  DFFPOSX1 arr_reg_0__23_ ( .D(n8325), .CLK(clk), .Q(arr[23]) );
  DFFPOSX1 arr_reg_0__22_ ( .D(n8324), .CLK(clk), .Q(arr[22]) );
  DFFPOSX1 arr_reg_0__21_ ( .D(n8323), .CLK(clk), .Q(arr[21]) );
  DFFPOSX1 arr_reg_0__20_ ( .D(n8322), .CLK(clk), .Q(arr[20]) );
  DFFPOSX1 arr_reg_0__19_ ( .D(n8321), .CLK(clk), .Q(arr[19]) );
  DFFPOSX1 arr_reg_0__18_ ( .D(n8320), .CLK(clk), .Q(arr[18]) );
  DFFPOSX1 arr_reg_0__17_ ( .D(n8319), .CLK(clk), .Q(arr[17]) );
  DFFPOSX1 arr_reg_0__16_ ( .D(n8318), .CLK(clk), .Q(arr[16]) );
  DFFPOSX1 arr_reg_0__15_ ( .D(n8317), .CLK(clk), .Q(arr[15]) );
  DFFPOSX1 arr_reg_0__14_ ( .D(n8316), .CLK(clk), .Q(arr[14]) );
  DFFPOSX1 arr_reg_0__13_ ( .D(n8315), .CLK(clk), .Q(arr[13]) );
  DFFPOSX1 arr_reg_0__12_ ( .D(n8314), .CLK(clk), .Q(arr[12]) );
  DFFPOSX1 arr_reg_0__11_ ( .D(n8313), .CLK(clk), .Q(arr[11]) );
  DFFPOSX1 arr_reg_0__10_ ( .D(n8312), .CLK(clk), .Q(arr[10]) );
  DFFPOSX1 arr_reg_0__9_ ( .D(n8311), .CLK(clk), .Q(arr[9]) );
  DFFPOSX1 arr_reg_0__8_ ( .D(n8310), .CLK(clk), .Q(arr[8]) );
  DFFPOSX1 arr_reg_0__7_ ( .D(n8309), .CLK(clk), .Q(arr[7]) );
  DFFPOSX1 arr_reg_0__6_ ( .D(n8308), .CLK(clk), .Q(arr[6]) );
  DFFPOSX1 arr_reg_0__5_ ( .D(n8307), .CLK(clk), .Q(arr[5]) );
  DFFPOSX1 arr_reg_0__4_ ( .D(n8306), .CLK(clk), .Q(arr[4]) );
  DFFPOSX1 arr_reg_0__3_ ( .D(n8305), .CLK(clk), .Q(arr[3]) );
  DFFPOSX1 arr_reg_0__2_ ( .D(n8304), .CLK(clk), .Q(arr[2]) );
  DFFPOSX1 arr_reg_0__1_ ( .D(n8303), .CLK(clk), .Q(arr[1]) );
  DFFPOSX1 arr_reg_0__0_ ( .D(n8302), .CLK(clk), .Q(arr[0]) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n8301), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n8300), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n8299), .CLK(clk), .Q(n15) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n8298), .CLK(clk), .Q(n16) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n8297), .CLK(clk), .Q(n17) );
  DFFPOSX1 rd_ptr_reg_5_ ( .D(n8296), .CLK(clk), .Q(n18) );
  AOI22X1 U4 ( .A(n2730), .B(n5482), .C(n3555), .D(n5483), .Y(n5481) );
  AOI22X1 U6 ( .A(n2729), .B(n5482), .C(n17), .D(n5483), .Y(n5484) );
  AOI22X1 U8 ( .A(n2728), .B(n5482), .C(n16), .D(n5483), .Y(n5485) );
  AOI22X1 U10 ( .A(n2727), .B(n5482), .C(n15), .D(n5483), .Y(n5486) );
  AOI22X1 U12 ( .A(n2726), .B(n5482), .C(n14), .D(n5483), .Y(n5487) );
  AOI22X1 U14 ( .A(n2725), .B(n5482), .C(n13), .D(n5483), .Y(n5488) );
  NOR2X1 U15 ( .A(n5483), .B(reset), .Y(n5482) );
  OAI21X1 U17 ( .A(n3549), .B(n5491), .C(n5492), .Y(n8302) );
  NAND2X1 U18 ( .A(arr[0]), .B(n3552), .Y(n5492) );
  OAI21X1 U19 ( .A(n3549), .B(n5493), .C(n5494), .Y(n8303) );
  NAND2X1 U20 ( .A(arr[1]), .B(n3552), .Y(n5494) );
  OAI21X1 U21 ( .A(n3549), .B(n5495), .C(n5496), .Y(n8304) );
  NAND2X1 U22 ( .A(arr[2]), .B(n3552), .Y(n5496) );
  OAI21X1 U23 ( .A(n3549), .B(n5497), .C(n5498), .Y(n8305) );
  NAND2X1 U24 ( .A(arr[3]), .B(n3552), .Y(n5498) );
  OAI21X1 U25 ( .A(n3549), .B(n5499), .C(n5500), .Y(n8306) );
  NAND2X1 U26 ( .A(arr[4]), .B(n3552), .Y(n5500) );
  OAI21X1 U27 ( .A(n3550), .B(n5501), .C(n5502), .Y(n8307) );
  NAND2X1 U28 ( .A(arr[5]), .B(n3552), .Y(n5502) );
  OAI21X1 U29 ( .A(n3550), .B(n5503), .C(n5504), .Y(n8308) );
  NAND2X1 U30 ( .A(arr[6]), .B(n3552), .Y(n5504) );
  OAI21X1 U31 ( .A(n3550), .B(n5505), .C(n5506), .Y(n8309) );
  NAND2X1 U32 ( .A(arr[7]), .B(n3552), .Y(n5506) );
  OAI21X1 U33 ( .A(n3549), .B(n5507), .C(n5508), .Y(n8310) );
  NAND2X1 U34 ( .A(arr[8]), .B(n3552), .Y(n5508) );
  OAI21X1 U35 ( .A(n3550), .B(n5509), .C(n5510), .Y(n8311) );
  NAND2X1 U36 ( .A(arr[9]), .B(n3552), .Y(n5510) );
  OAI21X1 U37 ( .A(n3551), .B(n5511), .C(n5512), .Y(n8312) );
  NAND2X1 U38 ( .A(arr[10]), .B(n3552), .Y(n5512) );
  OAI21X1 U39 ( .A(n3551), .B(n5513), .C(n5514), .Y(n8313) );
  NAND2X1 U40 ( .A(arr[11]), .B(n3552), .Y(n5514) );
  OAI21X1 U41 ( .A(n3551), .B(n5515), .C(n5516), .Y(n8314) );
  NAND2X1 U42 ( .A(arr[12]), .B(n3552), .Y(n5516) );
  OAI21X1 U43 ( .A(n3550), .B(n5517), .C(n5518), .Y(n8315) );
  NAND2X1 U44 ( .A(arr[13]), .B(n3553), .Y(n5518) );
  OAI21X1 U45 ( .A(n3552), .B(n5519), .C(n5520), .Y(n8316) );
  NAND2X1 U46 ( .A(arr[14]), .B(n3553), .Y(n5520) );
  OAI21X1 U47 ( .A(n3552), .B(n5521), .C(n5522), .Y(n8317) );
  NAND2X1 U48 ( .A(arr[15]), .B(n3553), .Y(n5522) );
  OAI21X1 U49 ( .A(n3551), .B(n5523), .C(n5524), .Y(n8318) );
  NAND2X1 U50 ( .A(arr[16]), .B(n3553), .Y(n5524) );
  OAI21X1 U51 ( .A(n3551), .B(n5525), .C(n5526), .Y(n8319) );
  NAND2X1 U52 ( .A(arr[17]), .B(n3553), .Y(n5526) );
  OAI21X1 U53 ( .A(n3551), .B(n5527), .C(n5528), .Y(n8320) );
  NAND2X1 U54 ( .A(arr[18]), .B(n3553), .Y(n5528) );
  OAI21X1 U55 ( .A(n3551), .B(n5529), .C(n5530), .Y(n8321) );
  NAND2X1 U56 ( .A(arr[19]), .B(n3553), .Y(n5530) );
  OAI21X1 U57 ( .A(n3551), .B(n5531), .C(n5532), .Y(n8322) );
  NAND2X1 U58 ( .A(arr[20]), .B(n3553), .Y(n5532) );
  OAI21X1 U59 ( .A(n3551), .B(n5533), .C(n5534), .Y(n8323) );
  NAND2X1 U60 ( .A(arr[21]), .B(n3553), .Y(n5534) );
  OAI21X1 U61 ( .A(n3551), .B(n5535), .C(n5536), .Y(n8324) );
  NAND2X1 U62 ( .A(arr[22]), .B(n3553), .Y(n5536) );
  OAI21X1 U63 ( .A(n3551), .B(n5537), .C(n5538), .Y(n8325) );
  NAND2X1 U64 ( .A(arr[23]), .B(n3553), .Y(n5538) );
  OAI21X1 U65 ( .A(n3551), .B(n5539), .C(n5540), .Y(n8326) );
  NAND2X1 U66 ( .A(arr[24]), .B(n3553), .Y(n5540) );
  OAI21X1 U67 ( .A(n3551), .B(n5541), .C(n5542), .Y(n8327) );
  NAND2X1 U68 ( .A(arr[25]), .B(n3553), .Y(n5542) );
  OAI21X1 U69 ( .A(n3550), .B(n5543), .C(n5544), .Y(n8328) );
  NAND2X1 U70 ( .A(arr[26]), .B(n3553), .Y(n5544) );
  OAI21X1 U71 ( .A(n3550), .B(n5545), .C(n5546), .Y(n8329) );
  NAND2X1 U72 ( .A(arr[27]), .B(n3553), .Y(n5546) );
  OAI21X1 U73 ( .A(n3550), .B(n5547), .C(n5548), .Y(n8330) );
  NAND2X1 U74 ( .A(arr[28]), .B(n3553), .Y(n5548) );
  OAI21X1 U75 ( .A(n3550), .B(n5549), .C(n5550), .Y(n8331) );
  NAND2X1 U76 ( .A(arr[29]), .B(n3554), .Y(n5550) );
  OAI21X1 U77 ( .A(n3550), .B(n5551), .C(n5552), .Y(n8332) );
  NAND2X1 U78 ( .A(arr[30]), .B(n3554), .Y(n5552) );
  OAI21X1 U79 ( .A(n3550), .B(n5553), .C(n5554), .Y(n8333) );
  NAND2X1 U80 ( .A(arr[31]), .B(n3554), .Y(n5554) );
  OAI21X1 U81 ( .A(n3550), .B(n5555), .C(n5556), .Y(n8334) );
  NAND2X1 U82 ( .A(arr[32]), .B(n3554), .Y(n5556) );
  OAI21X1 U83 ( .A(n3550), .B(n5557), .C(n5558), .Y(n8335) );
  NAND2X1 U84 ( .A(arr[33]), .B(n3554), .Y(n5558) );
  OAI21X1 U85 ( .A(n3549), .B(n5559), .C(n5560), .Y(n8336) );
  NAND2X1 U86 ( .A(arr[34]), .B(n3554), .Y(n5560) );
  OAI21X1 U87 ( .A(n3549), .B(n5561), .C(n5562), .Y(n8337) );
  NAND2X1 U88 ( .A(arr[35]), .B(n3554), .Y(n5562) );
  OAI21X1 U89 ( .A(n3549), .B(n5563), .C(n5564), .Y(n8338) );
  NAND2X1 U90 ( .A(arr[36]), .B(n3554), .Y(n5564) );
  OAI21X1 U91 ( .A(n3549), .B(n5565), .C(n5566), .Y(n8339) );
  NAND2X1 U92 ( .A(arr[37]), .B(n3554), .Y(n5566) );
  OAI21X1 U93 ( .A(n3549), .B(n5567), .C(n5568), .Y(n8340) );
  NAND2X1 U94 ( .A(arr[38]), .B(n3554), .Y(n5568) );
  OAI21X1 U95 ( .A(n3549), .B(n5569), .C(n5570), .Y(n8341) );
  NAND2X1 U96 ( .A(arr[39]), .B(n3552), .Y(n5570) );
  OAI21X1 U97 ( .A(n3549), .B(n5571), .C(n5572), .Y(n8342) );
  NAND2X1 U98 ( .A(arr[40]), .B(n3553), .Y(n5572) );
  NAND2X1 U99 ( .A(n5573), .B(n5574), .Y(n5490) );
  OAI21X1 U100 ( .A(n5491), .B(n3543), .C(n5576), .Y(n8343) );
  NAND2X1 U101 ( .A(arr[41]), .B(n3546), .Y(n5576) );
  OAI21X1 U102 ( .A(n5493), .B(n3543), .C(n5577), .Y(n8344) );
  NAND2X1 U103 ( .A(arr[42]), .B(n3546), .Y(n5577) );
  OAI21X1 U104 ( .A(n5495), .B(n3543), .C(n5578), .Y(n8345) );
  NAND2X1 U105 ( .A(arr[43]), .B(n3546), .Y(n5578) );
  OAI21X1 U106 ( .A(n5497), .B(n3543), .C(n5579), .Y(n8346) );
  NAND2X1 U107 ( .A(arr[44]), .B(n3546), .Y(n5579) );
  OAI21X1 U108 ( .A(n5499), .B(n3543), .C(n5580), .Y(n8347) );
  NAND2X1 U109 ( .A(arr[45]), .B(n3546), .Y(n5580) );
  OAI21X1 U110 ( .A(n5501), .B(n3544), .C(n5581), .Y(n8348) );
  NAND2X1 U111 ( .A(arr[46]), .B(n3546), .Y(n5581) );
  OAI21X1 U112 ( .A(n5503), .B(n3544), .C(n5582), .Y(n8349) );
  NAND2X1 U113 ( .A(arr[47]), .B(n3546), .Y(n5582) );
  OAI21X1 U114 ( .A(n5505), .B(n3544), .C(n5583), .Y(n8350) );
  NAND2X1 U115 ( .A(arr[48]), .B(n3546), .Y(n5583) );
  OAI21X1 U116 ( .A(n5507), .B(n3543), .C(n5584), .Y(n8351) );
  NAND2X1 U117 ( .A(arr[49]), .B(n3546), .Y(n5584) );
  OAI21X1 U118 ( .A(n5509), .B(n3544), .C(n5585), .Y(n8352) );
  NAND2X1 U119 ( .A(arr[50]), .B(n3546), .Y(n5585) );
  OAI21X1 U120 ( .A(n5511), .B(n3545), .C(n5586), .Y(n8353) );
  NAND2X1 U121 ( .A(arr[51]), .B(n3546), .Y(n5586) );
  OAI21X1 U122 ( .A(n5513), .B(n3545), .C(n5587), .Y(n8354) );
  NAND2X1 U123 ( .A(arr[52]), .B(n3546), .Y(n5587) );
  OAI21X1 U124 ( .A(n5515), .B(n3545), .C(n5588), .Y(n8355) );
  NAND2X1 U125 ( .A(arr[53]), .B(n3546), .Y(n5588) );
  OAI21X1 U126 ( .A(n5517), .B(n3544), .C(n5589), .Y(n8356) );
  NAND2X1 U127 ( .A(arr[54]), .B(n3547), .Y(n5589) );
  OAI21X1 U128 ( .A(n5519), .B(n3546), .C(n5590), .Y(n8357) );
  NAND2X1 U129 ( .A(arr[55]), .B(n3547), .Y(n5590) );
  OAI21X1 U130 ( .A(n5521), .B(n3546), .C(n5591), .Y(n8358) );
  NAND2X1 U131 ( .A(arr[56]), .B(n3547), .Y(n5591) );
  OAI21X1 U132 ( .A(n5523), .B(n3545), .C(n5592), .Y(n8359) );
  NAND2X1 U133 ( .A(arr[57]), .B(n3547), .Y(n5592) );
  OAI21X1 U134 ( .A(n5525), .B(n3545), .C(n5593), .Y(n8360) );
  NAND2X1 U135 ( .A(arr[58]), .B(n3547), .Y(n5593) );
  OAI21X1 U136 ( .A(n5527), .B(n3545), .C(n5594), .Y(n8361) );
  NAND2X1 U137 ( .A(arr[59]), .B(n3547), .Y(n5594) );
  OAI21X1 U138 ( .A(n5529), .B(n3545), .C(n5595), .Y(n8362) );
  NAND2X1 U139 ( .A(arr[60]), .B(n3547), .Y(n5595) );
  OAI21X1 U140 ( .A(n5531), .B(n3545), .C(n5596), .Y(n8363) );
  NAND2X1 U141 ( .A(arr[61]), .B(n3547), .Y(n5596) );
  OAI21X1 U142 ( .A(n5533), .B(n3545), .C(n5597), .Y(n8364) );
  NAND2X1 U143 ( .A(arr[62]), .B(n3547), .Y(n5597) );
  OAI21X1 U144 ( .A(n5535), .B(n3545), .C(n5598), .Y(n8365) );
  NAND2X1 U145 ( .A(arr[63]), .B(n3547), .Y(n5598) );
  OAI21X1 U146 ( .A(n5537), .B(n3545), .C(n5599), .Y(n8366) );
  NAND2X1 U147 ( .A(arr[64]), .B(n3547), .Y(n5599) );
  OAI21X1 U148 ( .A(n5539), .B(n3545), .C(n5600), .Y(n8367) );
  NAND2X1 U149 ( .A(arr[65]), .B(n3547), .Y(n5600) );
  OAI21X1 U150 ( .A(n5541), .B(n3545), .C(n5601), .Y(n8368) );
  NAND2X1 U151 ( .A(arr[66]), .B(n3547), .Y(n5601) );
  OAI21X1 U152 ( .A(n5543), .B(n3544), .C(n5602), .Y(n8369) );
  NAND2X1 U153 ( .A(arr[67]), .B(n3547), .Y(n5602) );
  OAI21X1 U154 ( .A(n5545), .B(n3544), .C(n5603), .Y(n8370) );
  NAND2X1 U155 ( .A(arr[68]), .B(n3547), .Y(n5603) );
  OAI21X1 U156 ( .A(n5547), .B(n3544), .C(n5604), .Y(n8371) );
  NAND2X1 U157 ( .A(arr[69]), .B(n3547), .Y(n5604) );
  OAI21X1 U158 ( .A(n5549), .B(n3544), .C(n5605), .Y(n8372) );
  NAND2X1 U159 ( .A(arr[70]), .B(n3547), .Y(n5605) );
  OAI21X1 U160 ( .A(n5551), .B(n3544), .C(n5606), .Y(n8373) );
  NAND2X1 U161 ( .A(arr[71]), .B(n3548), .Y(n5606) );
  OAI21X1 U162 ( .A(n5553), .B(n3544), .C(n5607), .Y(n8374) );
  NAND2X1 U163 ( .A(arr[72]), .B(n3548), .Y(n5607) );
  OAI21X1 U164 ( .A(n5555), .B(n3544), .C(n5608), .Y(n8375) );
  NAND2X1 U165 ( .A(arr[73]), .B(n3548), .Y(n5608) );
  OAI21X1 U166 ( .A(n5557), .B(n3544), .C(n5609), .Y(n8376) );
  NAND2X1 U167 ( .A(arr[74]), .B(n3548), .Y(n5609) );
  OAI21X1 U168 ( .A(n5559), .B(n3543), .C(n5610), .Y(n8377) );
  NAND2X1 U169 ( .A(arr[75]), .B(n3548), .Y(n5610) );
  OAI21X1 U170 ( .A(n5561), .B(n3543), .C(n5611), .Y(n8378) );
  NAND2X1 U171 ( .A(arr[76]), .B(n3548), .Y(n5611) );
  OAI21X1 U172 ( .A(n5563), .B(n3543), .C(n5612), .Y(n8379) );
  NAND2X1 U173 ( .A(arr[77]), .B(n3548), .Y(n5612) );
  OAI21X1 U174 ( .A(n5565), .B(n3543), .C(n5613), .Y(n8380) );
  NAND2X1 U175 ( .A(arr[78]), .B(n3548), .Y(n5613) );
  OAI21X1 U176 ( .A(n5567), .B(n3543), .C(n5614), .Y(n8381) );
  NAND2X1 U177 ( .A(arr[79]), .B(n3548), .Y(n5614) );
  OAI21X1 U178 ( .A(n5569), .B(n3543), .C(n5615), .Y(n8382) );
  NAND2X1 U179 ( .A(arr[80]), .B(n3546), .Y(n5615) );
  OAI21X1 U180 ( .A(n5571), .B(n3543), .C(n5616), .Y(n8383) );
  NAND2X1 U181 ( .A(arr[81]), .B(n3546), .Y(n5616) );
  NAND2X1 U182 ( .A(n5617), .B(n5574), .Y(n5575) );
  OAI21X1 U183 ( .A(n5491), .B(n3537), .C(n5619), .Y(n8384) );
  NAND2X1 U184 ( .A(arr[82]), .B(n3540), .Y(n5619) );
  OAI21X1 U185 ( .A(n5493), .B(n3537), .C(n5620), .Y(n8385) );
  NAND2X1 U186 ( .A(arr[83]), .B(n3540), .Y(n5620) );
  OAI21X1 U187 ( .A(n5495), .B(n3537), .C(n5621), .Y(n8386) );
  NAND2X1 U188 ( .A(arr[84]), .B(n3540), .Y(n5621) );
  OAI21X1 U189 ( .A(n5497), .B(n3537), .C(n5622), .Y(n8387) );
  NAND2X1 U190 ( .A(arr[85]), .B(n3540), .Y(n5622) );
  OAI21X1 U191 ( .A(n5499), .B(n3537), .C(n5623), .Y(n8388) );
  NAND2X1 U192 ( .A(arr[86]), .B(n3540), .Y(n5623) );
  OAI21X1 U193 ( .A(n5501), .B(n3538), .C(n5624), .Y(n8389) );
  NAND2X1 U194 ( .A(arr[87]), .B(n3540), .Y(n5624) );
  OAI21X1 U195 ( .A(n5503), .B(n3538), .C(n5625), .Y(n8390) );
  NAND2X1 U196 ( .A(arr[88]), .B(n3540), .Y(n5625) );
  OAI21X1 U197 ( .A(n5505), .B(n3538), .C(n5626), .Y(n8391) );
  NAND2X1 U198 ( .A(arr[89]), .B(n3540), .Y(n5626) );
  OAI21X1 U199 ( .A(n5507), .B(n3537), .C(n5627), .Y(n8392) );
  NAND2X1 U200 ( .A(arr[90]), .B(n3540), .Y(n5627) );
  OAI21X1 U201 ( .A(n5509), .B(n3538), .C(n5628), .Y(n8393) );
  NAND2X1 U202 ( .A(arr[91]), .B(n3540), .Y(n5628) );
  OAI21X1 U203 ( .A(n5511), .B(n3539), .C(n5629), .Y(n8394) );
  NAND2X1 U204 ( .A(arr[92]), .B(n3540), .Y(n5629) );
  OAI21X1 U205 ( .A(n5513), .B(n3539), .C(n5630), .Y(n8395) );
  NAND2X1 U206 ( .A(arr[93]), .B(n3540), .Y(n5630) );
  OAI21X1 U207 ( .A(n5515), .B(n3539), .C(n5631), .Y(n8396) );
  NAND2X1 U208 ( .A(arr[94]), .B(n3540), .Y(n5631) );
  OAI21X1 U209 ( .A(n5517), .B(n3538), .C(n5632), .Y(n8397) );
  NAND2X1 U210 ( .A(arr[95]), .B(n3541), .Y(n5632) );
  OAI21X1 U211 ( .A(n5519), .B(n3540), .C(n5633), .Y(n8398) );
  NAND2X1 U212 ( .A(arr[96]), .B(n3541), .Y(n5633) );
  OAI21X1 U213 ( .A(n5521), .B(n3540), .C(n5634), .Y(n8399) );
  NAND2X1 U214 ( .A(arr[97]), .B(n3541), .Y(n5634) );
  OAI21X1 U215 ( .A(n5523), .B(n3539), .C(n5635), .Y(n8400) );
  NAND2X1 U216 ( .A(arr[98]), .B(n3541), .Y(n5635) );
  OAI21X1 U217 ( .A(n5525), .B(n3539), .C(n5636), .Y(n8401) );
  NAND2X1 U218 ( .A(arr[99]), .B(n3541), .Y(n5636) );
  OAI21X1 U219 ( .A(n5527), .B(n3539), .C(n5637), .Y(n8402) );
  NAND2X1 U220 ( .A(arr[100]), .B(n3541), .Y(n5637) );
  OAI21X1 U221 ( .A(n5529), .B(n3539), .C(n5638), .Y(n8403) );
  NAND2X1 U222 ( .A(arr[101]), .B(n3541), .Y(n5638) );
  OAI21X1 U223 ( .A(n5531), .B(n3539), .C(n5639), .Y(n8404) );
  NAND2X1 U224 ( .A(arr[102]), .B(n3541), .Y(n5639) );
  OAI21X1 U225 ( .A(n5533), .B(n3539), .C(n5640), .Y(n8405) );
  NAND2X1 U226 ( .A(arr[103]), .B(n3541), .Y(n5640) );
  OAI21X1 U227 ( .A(n5535), .B(n3539), .C(n5641), .Y(n8406) );
  NAND2X1 U228 ( .A(arr[104]), .B(n3541), .Y(n5641) );
  OAI21X1 U229 ( .A(n5537), .B(n3539), .C(n5642), .Y(n8407) );
  NAND2X1 U230 ( .A(arr[105]), .B(n3541), .Y(n5642) );
  OAI21X1 U231 ( .A(n5539), .B(n3539), .C(n5643), .Y(n8408) );
  NAND2X1 U232 ( .A(arr[106]), .B(n3541), .Y(n5643) );
  OAI21X1 U233 ( .A(n5541), .B(n3539), .C(n5644), .Y(n8409) );
  NAND2X1 U234 ( .A(arr[107]), .B(n3541), .Y(n5644) );
  OAI21X1 U235 ( .A(n5543), .B(n3538), .C(n5645), .Y(n8410) );
  NAND2X1 U236 ( .A(arr[108]), .B(n3541), .Y(n5645) );
  OAI21X1 U237 ( .A(n5545), .B(n3538), .C(n5646), .Y(n8411) );
  NAND2X1 U238 ( .A(arr[109]), .B(n3541), .Y(n5646) );
  OAI21X1 U239 ( .A(n5547), .B(n3538), .C(n5647), .Y(n8412) );
  NAND2X1 U240 ( .A(arr[110]), .B(n3541), .Y(n5647) );
  OAI21X1 U241 ( .A(n5549), .B(n3538), .C(n5648), .Y(n8413) );
  NAND2X1 U242 ( .A(arr[111]), .B(n3541), .Y(n5648) );
  OAI21X1 U243 ( .A(n5551), .B(n3538), .C(n5649), .Y(n8414) );
  NAND2X1 U244 ( .A(arr[112]), .B(n3542), .Y(n5649) );
  OAI21X1 U245 ( .A(n5553), .B(n3538), .C(n5650), .Y(n8415) );
  NAND2X1 U246 ( .A(arr[113]), .B(n3542), .Y(n5650) );
  OAI21X1 U247 ( .A(n5555), .B(n3538), .C(n5651), .Y(n8416) );
  NAND2X1 U248 ( .A(arr[114]), .B(n3542), .Y(n5651) );
  OAI21X1 U249 ( .A(n5557), .B(n3538), .C(n5652), .Y(n8417) );
  NAND2X1 U250 ( .A(arr[115]), .B(n3542), .Y(n5652) );
  OAI21X1 U251 ( .A(n5559), .B(n3537), .C(n5653), .Y(n8418) );
  NAND2X1 U252 ( .A(arr[116]), .B(n3542), .Y(n5653) );
  OAI21X1 U253 ( .A(n5561), .B(n3537), .C(n5654), .Y(n8419) );
  NAND2X1 U254 ( .A(arr[117]), .B(n3542), .Y(n5654) );
  OAI21X1 U255 ( .A(n5563), .B(n3537), .C(n5655), .Y(n8420) );
  NAND2X1 U256 ( .A(arr[118]), .B(n3542), .Y(n5655) );
  OAI21X1 U257 ( .A(n5565), .B(n3537), .C(n5656), .Y(n8421) );
  NAND2X1 U258 ( .A(arr[119]), .B(n3542), .Y(n5656) );
  OAI21X1 U259 ( .A(n5567), .B(n3537), .C(n5657), .Y(n8422) );
  NAND2X1 U260 ( .A(arr[120]), .B(n3542), .Y(n5657) );
  OAI21X1 U261 ( .A(n5569), .B(n3537), .C(n5658), .Y(n8423) );
  NAND2X1 U262 ( .A(arr[121]), .B(n3540), .Y(n5658) );
  OAI21X1 U263 ( .A(n5571), .B(n3537), .C(n5659), .Y(n8424) );
  NAND2X1 U264 ( .A(arr[122]), .B(n3540), .Y(n5659) );
  NAND2X1 U265 ( .A(n5660), .B(n5574), .Y(n5618) );
  OAI21X1 U266 ( .A(n5491), .B(n3531), .C(n5662), .Y(n8425) );
  NAND2X1 U267 ( .A(arr[123]), .B(n3534), .Y(n5662) );
  OAI21X1 U268 ( .A(n5493), .B(n3531), .C(n5663), .Y(n8426) );
  NAND2X1 U269 ( .A(arr[124]), .B(n3534), .Y(n5663) );
  OAI21X1 U270 ( .A(n5495), .B(n3531), .C(n5664), .Y(n8427) );
  NAND2X1 U271 ( .A(arr[125]), .B(n3534), .Y(n5664) );
  OAI21X1 U272 ( .A(n5497), .B(n3531), .C(n5665), .Y(n8428) );
  NAND2X1 U273 ( .A(arr[126]), .B(n3534), .Y(n5665) );
  OAI21X1 U274 ( .A(n5499), .B(n3531), .C(n5666), .Y(n8429) );
  NAND2X1 U275 ( .A(arr[127]), .B(n3534), .Y(n5666) );
  OAI21X1 U276 ( .A(n5501), .B(n3532), .C(n5667), .Y(n8430) );
  NAND2X1 U277 ( .A(arr[128]), .B(n3534), .Y(n5667) );
  OAI21X1 U278 ( .A(n5503), .B(n3532), .C(n5668), .Y(n8431) );
  NAND2X1 U279 ( .A(arr[129]), .B(n3534), .Y(n5668) );
  OAI21X1 U280 ( .A(n5505), .B(n3532), .C(n5669), .Y(n8432) );
  NAND2X1 U281 ( .A(arr[130]), .B(n3534), .Y(n5669) );
  OAI21X1 U282 ( .A(n5507), .B(n3531), .C(n5670), .Y(n8433) );
  NAND2X1 U283 ( .A(arr[131]), .B(n3534), .Y(n5670) );
  OAI21X1 U284 ( .A(n5509), .B(n3532), .C(n5671), .Y(n8434) );
  NAND2X1 U285 ( .A(arr[132]), .B(n3534), .Y(n5671) );
  OAI21X1 U286 ( .A(n5511), .B(n3533), .C(n5672), .Y(n8435) );
  NAND2X1 U287 ( .A(arr[133]), .B(n3534), .Y(n5672) );
  OAI21X1 U288 ( .A(n5513), .B(n3533), .C(n5673), .Y(n8436) );
  NAND2X1 U289 ( .A(arr[134]), .B(n3534), .Y(n5673) );
  OAI21X1 U290 ( .A(n5515), .B(n3533), .C(n5674), .Y(n8437) );
  NAND2X1 U291 ( .A(arr[135]), .B(n3534), .Y(n5674) );
  OAI21X1 U292 ( .A(n5517), .B(n3532), .C(n5675), .Y(n8438) );
  NAND2X1 U293 ( .A(arr[136]), .B(n3535), .Y(n5675) );
  OAI21X1 U294 ( .A(n5519), .B(n3534), .C(n5676), .Y(n8439) );
  NAND2X1 U295 ( .A(arr[137]), .B(n3535), .Y(n5676) );
  OAI21X1 U296 ( .A(n5521), .B(n3534), .C(n5677), .Y(n8440) );
  NAND2X1 U297 ( .A(arr[138]), .B(n3535), .Y(n5677) );
  OAI21X1 U298 ( .A(n5523), .B(n3533), .C(n5678), .Y(n8441) );
  NAND2X1 U299 ( .A(arr[139]), .B(n3535), .Y(n5678) );
  OAI21X1 U300 ( .A(n5525), .B(n3533), .C(n5679), .Y(n8442) );
  NAND2X1 U301 ( .A(arr[140]), .B(n3535), .Y(n5679) );
  OAI21X1 U302 ( .A(n5527), .B(n3533), .C(n5680), .Y(n8443) );
  NAND2X1 U303 ( .A(arr[141]), .B(n3535), .Y(n5680) );
  OAI21X1 U304 ( .A(n5529), .B(n3533), .C(n5681), .Y(n8444) );
  NAND2X1 U305 ( .A(arr[142]), .B(n3535), .Y(n5681) );
  OAI21X1 U306 ( .A(n5531), .B(n3533), .C(n5682), .Y(n8445) );
  NAND2X1 U307 ( .A(arr[143]), .B(n3535), .Y(n5682) );
  OAI21X1 U308 ( .A(n5533), .B(n3533), .C(n5683), .Y(n8446) );
  NAND2X1 U309 ( .A(arr[144]), .B(n3535), .Y(n5683) );
  OAI21X1 U310 ( .A(n5535), .B(n3533), .C(n5684), .Y(n8447) );
  NAND2X1 U311 ( .A(arr[145]), .B(n3535), .Y(n5684) );
  OAI21X1 U312 ( .A(n5537), .B(n3533), .C(n5685), .Y(n8448) );
  NAND2X1 U313 ( .A(arr[146]), .B(n3535), .Y(n5685) );
  OAI21X1 U314 ( .A(n5539), .B(n3533), .C(n5686), .Y(n8449) );
  NAND2X1 U315 ( .A(arr[147]), .B(n3535), .Y(n5686) );
  OAI21X1 U316 ( .A(n5541), .B(n3533), .C(n5687), .Y(n8450) );
  NAND2X1 U317 ( .A(arr[148]), .B(n3535), .Y(n5687) );
  OAI21X1 U318 ( .A(n5543), .B(n3532), .C(n5688), .Y(n8451) );
  NAND2X1 U319 ( .A(arr[149]), .B(n3535), .Y(n5688) );
  OAI21X1 U320 ( .A(n5545), .B(n3532), .C(n5689), .Y(n8452) );
  NAND2X1 U321 ( .A(arr[150]), .B(n3535), .Y(n5689) );
  OAI21X1 U322 ( .A(n5547), .B(n3532), .C(n5690), .Y(n8453) );
  NAND2X1 U323 ( .A(arr[151]), .B(n3535), .Y(n5690) );
  OAI21X1 U324 ( .A(n5549), .B(n3532), .C(n5691), .Y(n8454) );
  NAND2X1 U325 ( .A(arr[152]), .B(n3535), .Y(n5691) );
  OAI21X1 U326 ( .A(n5551), .B(n3532), .C(n5692), .Y(n8455) );
  NAND2X1 U327 ( .A(arr[153]), .B(n3536), .Y(n5692) );
  OAI21X1 U328 ( .A(n5553), .B(n3532), .C(n5693), .Y(n8456) );
  NAND2X1 U329 ( .A(arr[154]), .B(n3536), .Y(n5693) );
  OAI21X1 U330 ( .A(n5555), .B(n3532), .C(n5694), .Y(n8457) );
  NAND2X1 U331 ( .A(arr[155]), .B(n3536), .Y(n5694) );
  OAI21X1 U332 ( .A(n5557), .B(n3532), .C(n5695), .Y(n8458) );
  NAND2X1 U333 ( .A(arr[156]), .B(n3536), .Y(n5695) );
  OAI21X1 U334 ( .A(n5559), .B(n3531), .C(n5696), .Y(n8459) );
  NAND2X1 U335 ( .A(arr[157]), .B(n3536), .Y(n5696) );
  OAI21X1 U336 ( .A(n5561), .B(n3531), .C(n5697), .Y(n8460) );
  NAND2X1 U337 ( .A(arr[158]), .B(n3536), .Y(n5697) );
  OAI21X1 U338 ( .A(n5563), .B(n3531), .C(n5698), .Y(n8461) );
  NAND2X1 U339 ( .A(arr[159]), .B(n3536), .Y(n5698) );
  OAI21X1 U340 ( .A(n5565), .B(n3531), .C(n5699), .Y(n8462) );
  NAND2X1 U341 ( .A(arr[160]), .B(n3536), .Y(n5699) );
  OAI21X1 U342 ( .A(n5567), .B(n3531), .C(n5700), .Y(n8463) );
  NAND2X1 U343 ( .A(arr[161]), .B(n3536), .Y(n5700) );
  OAI21X1 U344 ( .A(n5569), .B(n3531), .C(n5701), .Y(n8464) );
  NAND2X1 U345 ( .A(arr[162]), .B(n3534), .Y(n5701) );
  OAI21X1 U346 ( .A(n5571), .B(n3531), .C(n5702), .Y(n8465) );
  NAND2X1 U347 ( .A(arr[163]), .B(n3534), .Y(n5702) );
  NAND2X1 U348 ( .A(n5703), .B(n5574), .Y(n5661) );
  OAI21X1 U350 ( .A(n5491), .B(n3525), .C(n5707), .Y(n8466) );
  NAND2X1 U351 ( .A(arr[164]), .B(n3528), .Y(n5707) );
  OAI21X1 U352 ( .A(n5493), .B(n3525), .C(n5708), .Y(n8467) );
  NAND2X1 U353 ( .A(arr[165]), .B(n3528), .Y(n5708) );
  OAI21X1 U354 ( .A(n5495), .B(n3525), .C(n5709), .Y(n8468) );
  NAND2X1 U355 ( .A(arr[166]), .B(n3528), .Y(n5709) );
  OAI21X1 U356 ( .A(n5497), .B(n3525), .C(n5710), .Y(n8469) );
  NAND2X1 U357 ( .A(arr[167]), .B(n3528), .Y(n5710) );
  OAI21X1 U358 ( .A(n5499), .B(n3525), .C(n5711), .Y(n8470) );
  NAND2X1 U359 ( .A(arr[168]), .B(n3528), .Y(n5711) );
  OAI21X1 U360 ( .A(n5501), .B(n3526), .C(n5712), .Y(n8471) );
  NAND2X1 U361 ( .A(arr[169]), .B(n3528), .Y(n5712) );
  OAI21X1 U362 ( .A(n5503), .B(n3526), .C(n5713), .Y(n8472) );
  NAND2X1 U363 ( .A(arr[170]), .B(n3528), .Y(n5713) );
  OAI21X1 U364 ( .A(n5505), .B(n3526), .C(n5714), .Y(n8473) );
  NAND2X1 U365 ( .A(arr[171]), .B(n3528), .Y(n5714) );
  OAI21X1 U366 ( .A(n5507), .B(n3525), .C(n5715), .Y(n8474) );
  NAND2X1 U367 ( .A(arr[172]), .B(n3528), .Y(n5715) );
  OAI21X1 U368 ( .A(n5509), .B(n3526), .C(n5716), .Y(n8475) );
  NAND2X1 U369 ( .A(arr[173]), .B(n3528), .Y(n5716) );
  OAI21X1 U370 ( .A(n5511), .B(n3527), .C(n5717), .Y(n8476) );
  NAND2X1 U371 ( .A(arr[174]), .B(n3528), .Y(n5717) );
  OAI21X1 U372 ( .A(n5513), .B(n3527), .C(n5718), .Y(n8477) );
  NAND2X1 U373 ( .A(arr[175]), .B(n3528), .Y(n5718) );
  OAI21X1 U374 ( .A(n5515), .B(n3527), .C(n5719), .Y(n8478) );
  NAND2X1 U375 ( .A(arr[176]), .B(n3528), .Y(n5719) );
  OAI21X1 U376 ( .A(n5517), .B(n3526), .C(n5720), .Y(n8479) );
  NAND2X1 U377 ( .A(arr[177]), .B(n3529), .Y(n5720) );
  OAI21X1 U378 ( .A(n5519), .B(n3528), .C(n5721), .Y(n8480) );
  NAND2X1 U379 ( .A(arr[178]), .B(n3529), .Y(n5721) );
  OAI21X1 U380 ( .A(n5521), .B(n3528), .C(n5722), .Y(n8481) );
  NAND2X1 U381 ( .A(arr[179]), .B(n3529), .Y(n5722) );
  OAI21X1 U382 ( .A(n5523), .B(n3527), .C(n5723), .Y(n8482) );
  NAND2X1 U383 ( .A(arr[180]), .B(n3529), .Y(n5723) );
  OAI21X1 U384 ( .A(n5525), .B(n3527), .C(n5724), .Y(n8483) );
  NAND2X1 U385 ( .A(arr[181]), .B(n3529), .Y(n5724) );
  OAI21X1 U386 ( .A(n5527), .B(n3527), .C(n5725), .Y(n8484) );
  NAND2X1 U387 ( .A(arr[182]), .B(n3529), .Y(n5725) );
  OAI21X1 U388 ( .A(n5529), .B(n3527), .C(n5726), .Y(n8485) );
  NAND2X1 U389 ( .A(arr[183]), .B(n3529), .Y(n5726) );
  OAI21X1 U390 ( .A(n5531), .B(n3527), .C(n5727), .Y(n8486) );
  NAND2X1 U391 ( .A(arr[184]), .B(n3529), .Y(n5727) );
  OAI21X1 U392 ( .A(n5533), .B(n3527), .C(n5728), .Y(n8487) );
  NAND2X1 U393 ( .A(arr[185]), .B(n3529), .Y(n5728) );
  OAI21X1 U394 ( .A(n5535), .B(n3527), .C(n5729), .Y(n8488) );
  NAND2X1 U395 ( .A(arr[186]), .B(n3529), .Y(n5729) );
  OAI21X1 U396 ( .A(n5537), .B(n3527), .C(n5730), .Y(n8489) );
  NAND2X1 U397 ( .A(arr[187]), .B(n3529), .Y(n5730) );
  OAI21X1 U398 ( .A(n5539), .B(n3527), .C(n5731), .Y(n8490) );
  NAND2X1 U399 ( .A(arr[188]), .B(n3529), .Y(n5731) );
  OAI21X1 U400 ( .A(n5541), .B(n3527), .C(n5732), .Y(n8491) );
  NAND2X1 U401 ( .A(arr[189]), .B(n3529), .Y(n5732) );
  OAI21X1 U402 ( .A(n5543), .B(n3526), .C(n5733), .Y(n8492) );
  NAND2X1 U403 ( .A(arr[190]), .B(n3529), .Y(n5733) );
  OAI21X1 U404 ( .A(n5545), .B(n3526), .C(n5734), .Y(n8493) );
  NAND2X1 U405 ( .A(arr[191]), .B(n3529), .Y(n5734) );
  OAI21X1 U406 ( .A(n5547), .B(n3526), .C(n5735), .Y(n8494) );
  NAND2X1 U407 ( .A(arr[192]), .B(n3529), .Y(n5735) );
  OAI21X1 U408 ( .A(n5549), .B(n3526), .C(n5736), .Y(n8495) );
  NAND2X1 U409 ( .A(arr[193]), .B(n3529), .Y(n5736) );
  OAI21X1 U410 ( .A(n5551), .B(n3526), .C(n5737), .Y(n8496) );
  NAND2X1 U411 ( .A(arr[194]), .B(n3530), .Y(n5737) );
  OAI21X1 U412 ( .A(n5553), .B(n3526), .C(n5738), .Y(n8497) );
  NAND2X1 U413 ( .A(arr[195]), .B(n3530), .Y(n5738) );
  OAI21X1 U414 ( .A(n5555), .B(n3526), .C(n5739), .Y(n8498) );
  NAND2X1 U415 ( .A(arr[196]), .B(n3530), .Y(n5739) );
  OAI21X1 U416 ( .A(n5557), .B(n3526), .C(n5740), .Y(n8499) );
  NAND2X1 U417 ( .A(arr[197]), .B(n3530), .Y(n5740) );
  OAI21X1 U418 ( .A(n5559), .B(n3525), .C(n5741), .Y(n8500) );
  NAND2X1 U419 ( .A(arr[198]), .B(n3530), .Y(n5741) );
  OAI21X1 U420 ( .A(n5561), .B(n3525), .C(n5742), .Y(n8501) );
  NAND2X1 U421 ( .A(arr[199]), .B(n3530), .Y(n5742) );
  OAI21X1 U422 ( .A(n5563), .B(n3525), .C(n5743), .Y(n8502) );
  NAND2X1 U423 ( .A(arr[200]), .B(n3530), .Y(n5743) );
  OAI21X1 U424 ( .A(n5565), .B(n3525), .C(n5744), .Y(n8503) );
  NAND2X1 U425 ( .A(arr[201]), .B(n3530), .Y(n5744) );
  OAI21X1 U426 ( .A(n5567), .B(n3525), .C(n5745), .Y(n8504) );
  NAND2X1 U427 ( .A(arr[202]), .B(n3530), .Y(n5745) );
  OAI21X1 U428 ( .A(n5569), .B(n3525), .C(n5746), .Y(n8505) );
  NAND2X1 U429 ( .A(arr[203]), .B(n3528), .Y(n5746) );
  OAI21X1 U430 ( .A(n5571), .B(n3525), .C(n5747), .Y(n8506) );
  NAND2X1 U431 ( .A(arr[204]), .B(n3528), .Y(n5747) );
  NAND2X1 U432 ( .A(n5748), .B(n5573), .Y(n5706) );
  OAI21X1 U433 ( .A(n5491), .B(n3519), .C(n5750), .Y(n8507) );
  NAND2X1 U434 ( .A(arr[205]), .B(n3522), .Y(n5750) );
  OAI21X1 U435 ( .A(n5493), .B(n3519), .C(n5751), .Y(n8508) );
  NAND2X1 U436 ( .A(arr[206]), .B(n3522), .Y(n5751) );
  OAI21X1 U437 ( .A(n5495), .B(n3519), .C(n5752), .Y(n8509) );
  NAND2X1 U438 ( .A(arr[207]), .B(n3522), .Y(n5752) );
  OAI21X1 U439 ( .A(n5497), .B(n3519), .C(n5753), .Y(n8510) );
  NAND2X1 U440 ( .A(arr[208]), .B(n3522), .Y(n5753) );
  OAI21X1 U441 ( .A(n5499), .B(n3519), .C(n5754), .Y(n8511) );
  NAND2X1 U442 ( .A(arr[209]), .B(n3522), .Y(n5754) );
  OAI21X1 U443 ( .A(n5501), .B(n3520), .C(n5755), .Y(n8512) );
  NAND2X1 U444 ( .A(arr[210]), .B(n3522), .Y(n5755) );
  OAI21X1 U445 ( .A(n5503), .B(n3520), .C(n5756), .Y(n8513) );
  NAND2X1 U446 ( .A(arr[211]), .B(n3522), .Y(n5756) );
  OAI21X1 U447 ( .A(n5505), .B(n3520), .C(n5757), .Y(n8514) );
  NAND2X1 U448 ( .A(arr[212]), .B(n3522), .Y(n5757) );
  OAI21X1 U449 ( .A(n5507), .B(n3519), .C(n5758), .Y(n8515) );
  NAND2X1 U450 ( .A(arr[213]), .B(n3522), .Y(n5758) );
  OAI21X1 U451 ( .A(n5509), .B(n3520), .C(n5759), .Y(n8516) );
  NAND2X1 U452 ( .A(arr[214]), .B(n3522), .Y(n5759) );
  OAI21X1 U453 ( .A(n5511), .B(n3521), .C(n5760), .Y(n8517) );
  NAND2X1 U454 ( .A(arr[215]), .B(n3522), .Y(n5760) );
  OAI21X1 U455 ( .A(n5513), .B(n3521), .C(n5761), .Y(n8518) );
  NAND2X1 U456 ( .A(arr[216]), .B(n3522), .Y(n5761) );
  OAI21X1 U457 ( .A(n5515), .B(n3521), .C(n5762), .Y(n8519) );
  NAND2X1 U458 ( .A(arr[217]), .B(n3522), .Y(n5762) );
  OAI21X1 U459 ( .A(n5517), .B(n3520), .C(n5763), .Y(n8520) );
  NAND2X1 U460 ( .A(arr[218]), .B(n3523), .Y(n5763) );
  OAI21X1 U461 ( .A(n5519), .B(n3522), .C(n5764), .Y(n8521) );
  NAND2X1 U462 ( .A(arr[219]), .B(n3523), .Y(n5764) );
  OAI21X1 U463 ( .A(n5521), .B(n3522), .C(n5765), .Y(n8522) );
  NAND2X1 U464 ( .A(arr[220]), .B(n3523), .Y(n5765) );
  OAI21X1 U465 ( .A(n5523), .B(n3521), .C(n5766), .Y(n8523) );
  NAND2X1 U466 ( .A(arr[221]), .B(n3523), .Y(n5766) );
  OAI21X1 U467 ( .A(n5525), .B(n3521), .C(n5767), .Y(n8524) );
  NAND2X1 U468 ( .A(arr[222]), .B(n3523), .Y(n5767) );
  OAI21X1 U469 ( .A(n5527), .B(n3521), .C(n5768), .Y(n8525) );
  NAND2X1 U470 ( .A(arr[223]), .B(n3523), .Y(n5768) );
  OAI21X1 U471 ( .A(n5529), .B(n3521), .C(n5769), .Y(n8526) );
  NAND2X1 U472 ( .A(arr[224]), .B(n3523), .Y(n5769) );
  OAI21X1 U473 ( .A(n5531), .B(n3521), .C(n5770), .Y(n8527) );
  NAND2X1 U474 ( .A(arr[225]), .B(n3523), .Y(n5770) );
  OAI21X1 U475 ( .A(n5533), .B(n3521), .C(n5771), .Y(n8528) );
  NAND2X1 U476 ( .A(arr[226]), .B(n3523), .Y(n5771) );
  OAI21X1 U477 ( .A(n5535), .B(n3521), .C(n5772), .Y(n8529) );
  NAND2X1 U478 ( .A(arr[227]), .B(n3523), .Y(n5772) );
  OAI21X1 U479 ( .A(n5537), .B(n3521), .C(n5773), .Y(n8530) );
  NAND2X1 U480 ( .A(arr[228]), .B(n3523), .Y(n5773) );
  OAI21X1 U481 ( .A(n5539), .B(n3521), .C(n5774), .Y(n8531) );
  NAND2X1 U482 ( .A(arr[229]), .B(n3523), .Y(n5774) );
  OAI21X1 U483 ( .A(n5541), .B(n3521), .C(n5775), .Y(n8532) );
  NAND2X1 U484 ( .A(arr[230]), .B(n3523), .Y(n5775) );
  OAI21X1 U485 ( .A(n5543), .B(n3520), .C(n5776), .Y(n8533) );
  NAND2X1 U486 ( .A(arr[231]), .B(n3523), .Y(n5776) );
  OAI21X1 U487 ( .A(n5545), .B(n3520), .C(n5777), .Y(n8534) );
  NAND2X1 U488 ( .A(arr[232]), .B(n3523), .Y(n5777) );
  OAI21X1 U489 ( .A(n5547), .B(n3520), .C(n5778), .Y(n8535) );
  NAND2X1 U490 ( .A(arr[233]), .B(n3523), .Y(n5778) );
  OAI21X1 U491 ( .A(n5549), .B(n3520), .C(n5779), .Y(n8536) );
  NAND2X1 U492 ( .A(arr[234]), .B(n3523), .Y(n5779) );
  OAI21X1 U493 ( .A(n5551), .B(n3520), .C(n5780), .Y(n8537) );
  NAND2X1 U494 ( .A(arr[235]), .B(n3524), .Y(n5780) );
  OAI21X1 U495 ( .A(n5553), .B(n3520), .C(n5781), .Y(n8538) );
  NAND2X1 U496 ( .A(arr[236]), .B(n3524), .Y(n5781) );
  OAI21X1 U497 ( .A(n5555), .B(n3520), .C(n5782), .Y(n8539) );
  NAND2X1 U498 ( .A(arr[237]), .B(n3524), .Y(n5782) );
  OAI21X1 U499 ( .A(n5557), .B(n3520), .C(n5783), .Y(n8540) );
  NAND2X1 U500 ( .A(arr[238]), .B(n3524), .Y(n5783) );
  OAI21X1 U501 ( .A(n5559), .B(n3519), .C(n5784), .Y(n8541) );
  NAND2X1 U502 ( .A(arr[239]), .B(n3524), .Y(n5784) );
  OAI21X1 U503 ( .A(n5561), .B(n3519), .C(n5785), .Y(n8542) );
  NAND2X1 U504 ( .A(arr[240]), .B(n3524), .Y(n5785) );
  OAI21X1 U505 ( .A(n5563), .B(n3519), .C(n5786), .Y(n8543) );
  NAND2X1 U506 ( .A(arr[241]), .B(n3524), .Y(n5786) );
  OAI21X1 U507 ( .A(n5565), .B(n3519), .C(n5787), .Y(n8544) );
  NAND2X1 U508 ( .A(arr[242]), .B(n3524), .Y(n5787) );
  OAI21X1 U509 ( .A(n5567), .B(n3519), .C(n5788), .Y(n8545) );
  NAND2X1 U510 ( .A(arr[243]), .B(n3524), .Y(n5788) );
  OAI21X1 U511 ( .A(n5569), .B(n3519), .C(n5789), .Y(n8546) );
  NAND2X1 U512 ( .A(arr[244]), .B(n3522), .Y(n5789) );
  OAI21X1 U513 ( .A(n5571), .B(n3519), .C(n5790), .Y(n8547) );
  NAND2X1 U514 ( .A(arr[245]), .B(n3522), .Y(n5790) );
  NAND2X1 U515 ( .A(n5748), .B(n5617), .Y(n5749) );
  OAI21X1 U516 ( .A(n5491), .B(n3513), .C(n5792), .Y(n8548) );
  NAND2X1 U517 ( .A(arr[246]), .B(n3516), .Y(n5792) );
  OAI21X1 U518 ( .A(n5493), .B(n3513), .C(n5793), .Y(n8549) );
  NAND2X1 U519 ( .A(arr[247]), .B(n3516), .Y(n5793) );
  OAI21X1 U520 ( .A(n5495), .B(n3513), .C(n5794), .Y(n8550) );
  NAND2X1 U521 ( .A(arr[248]), .B(n3516), .Y(n5794) );
  OAI21X1 U522 ( .A(n5497), .B(n3513), .C(n5795), .Y(n8551) );
  NAND2X1 U523 ( .A(arr[249]), .B(n3516), .Y(n5795) );
  OAI21X1 U524 ( .A(n5499), .B(n3513), .C(n5796), .Y(n8552) );
  NAND2X1 U525 ( .A(arr[250]), .B(n3516), .Y(n5796) );
  OAI21X1 U526 ( .A(n5501), .B(n3514), .C(n5797), .Y(n8553) );
  NAND2X1 U527 ( .A(arr[251]), .B(n3516), .Y(n5797) );
  OAI21X1 U528 ( .A(n5503), .B(n3514), .C(n5798), .Y(n8554) );
  NAND2X1 U529 ( .A(arr[252]), .B(n3516), .Y(n5798) );
  OAI21X1 U530 ( .A(n5505), .B(n3514), .C(n5799), .Y(n8555) );
  NAND2X1 U531 ( .A(arr[253]), .B(n3516), .Y(n5799) );
  OAI21X1 U532 ( .A(n5507), .B(n3513), .C(n5800), .Y(n8556) );
  NAND2X1 U533 ( .A(arr[254]), .B(n3516), .Y(n5800) );
  OAI21X1 U534 ( .A(n5509), .B(n3514), .C(n5801), .Y(n8557) );
  NAND2X1 U535 ( .A(arr[255]), .B(n3516), .Y(n5801) );
  OAI21X1 U536 ( .A(n5511), .B(n3515), .C(n5802), .Y(n8558) );
  NAND2X1 U537 ( .A(arr[256]), .B(n3516), .Y(n5802) );
  OAI21X1 U538 ( .A(n5513), .B(n3515), .C(n5803), .Y(n8559) );
  NAND2X1 U539 ( .A(arr[257]), .B(n3516), .Y(n5803) );
  OAI21X1 U540 ( .A(n5515), .B(n3515), .C(n5804), .Y(n8560) );
  NAND2X1 U541 ( .A(arr[258]), .B(n3516), .Y(n5804) );
  OAI21X1 U542 ( .A(n5517), .B(n3514), .C(n5805), .Y(n8561) );
  NAND2X1 U543 ( .A(arr[259]), .B(n3517), .Y(n5805) );
  OAI21X1 U544 ( .A(n5519), .B(n3516), .C(n5806), .Y(n8562) );
  NAND2X1 U545 ( .A(arr[260]), .B(n3517), .Y(n5806) );
  OAI21X1 U546 ( .A(n5521), .B(n3516), .C(n5807), .Y(n8563) );
  NAND2X1 U547 ( .A(arr[261]), .B(n3517), .Y(n5807) );
  OAI21X1 U548 ( .A(n5523), .B(n3515), .C(n5808), .Y(n8564) );
  NAND2X1 U549 ( .A(arr[262]), .B(n3517), .Y(n5808) );
  OAI21X1 U550 ( .A(n5525), .B(n3515), .C(n5809), .Y(n8565) );
  NAND2X1 U551 ( .A(arr[263]), .B(n3517), .Y(n5809) );
  OAI21X1 U552 ( .A(n5527), .B(n3515), .C(n5810), .Y(n8566) );
  NAND2X1 U553 ( .A(arr[264]), .B(n3517), .Y(n5810) );
  OAI21X1 U554 ( .A(n5529), .B(n3515), .C(n5811), .Y(n8567) );
  NAND2X1 U555 ( .A(arr[265]), .B(n3517), .Y(n5811) );
  OAI21X1 U556 ( .A(n5531), .B(n3515), .C(n5812), .Y(n8568) );
  NAND2X1 U557 ( .A(arr[266]), .B(n3517), .Y(n5812) );
  OAI21X1 U558 ( .A(n5533), .B(n3515), .C(n5813), .Y(n8569) );
  NAND2X1 U559 ( .A(arr[267]), .B(n3517), .Y(n5813) );
  OAI21X1 U560 ( .A(n5535), .B(n3515), .C(n5814), .Y(n8570) );
  NAND2X1 U561 ( .A(arr[268]), .B(n3517), .Y(n5814) );
  OAI21X1 U562 ( .A(n5537), .B(n3515), .C(n5815), .Y(n8571) );
  NAND2X1 U563 ( .A(arr[269]), .B(n3517), .Y(n5815) );
  OAI21X1 U564 ( .A(n5539), .B(n3515), .C(n5816), .Y(n8572) );
  NAND2X1 U565 ( .A(arr[270]), .B(n3517), .Y(n5816) );
  OAI21X1 U566 ( .A(n5541), .B(n3515), .C(n5817), .Y(n8573) );
  NAND2X1 U567 ( .A(arr[271]), .B(n3517), .Y(n5817) );
  OAI21X1 U568 ( .A(n5543), .B(n3514), .C(n5818), .Y(n8574) );
  NAND2X1 U569 ( .A(arr[272]), .B(n3517), .Y(n5818) );
  OAI21X1 U570 ( .A(n5545), .B(n3514), .C(n5819), .Y(n8575) );
  NAND2X1 U571 ( .A(arr[273]), .B(n3517), .Y(n5819) );
  OAI21X1 U572 ( .A(n5547), .B(n3514), .C(n5820), .Y(n8576) );
  NAND2X1 U573 ( .A(arr[274]), .B(n3517), .Y(n5820) );
  OAI21X1 U574 ( .A(n5549), .B(n3514), .C(n5821), .Y(n8577) );
  NAND2X1 U575 ( .A(arr[275]), .B(n3517), .Y(n5821) );
  OAI21X1 U576 ( .A(n5551), .B(n3514), .C(n5822), .Y(n8578) );
  NAND2X1 U577 ( .A(arr[276]), .B(n3518), .Y(n5822) );
  OAI21X1 U578 ( .A(n5553), .B(n3514), .C(n5823), .Y(n8579) );
  NAND2X1 U579 ( .A(arr[277]), .B(n3518), .Y(n5823) );
  OAI21X1 U580 ( .A(n5555), .B(n3514), .C(n5824), .Y(n8580) );
  NAND2X1 U581 ( .A(arr[278]), .B(n3518), .Y(n5824) );
  OAI21X1 U582 ( .A(n5557), .B(n3514), .C(n5825), .Y(n8581) );
  NAND2X1 U583 ( .A(arr[279]), .B(n3518), .Y(n5825) );
  OAI21X1 U584 ( .A(n5559), .B(n3513), .C(n5826), .Y(n8582) );
  NAND2X1 U585 ( .A(arr[280]), .B(n3518), .Y(n5826) );
  OAI21X1 U586 ( .A(n5561), .B(n3513), .C(n5827), .Y(n8583) );
  NAND2X1 U587 ( .A(arr[281]), .B(n3518), .Y(n5827) );
  OAI21X1 U588 ( .A(n5563), .B(n3513), .C(n5828), .Y(n8584) );
  NAND2X1 U589 ( .A(arr[282]), .B(n3518), .Y(n5828) );
  OAI21X1 U590 ( .A(n5565), .B(n3513), .C(n5829), .Y(n8585) );
  NAND2X1 U591 ( .A(arr[283]), .B(n3518), .Y(n5829) );
  OAI21X1 U592 ( .A(n5567), .B(n3513), .C(n5830), .Y(n8586) );
  NAND2X1 U593 ( .A(arr[284]), .B(n3518), .Y(n5830) );
  OAI21X1 U594 ( .A(n5569), .B(n3513), .C(n5831), .Y(n8587) );
  NAND2X1 U595 ( .A(arr[285]), .B(n3516), .Y(n5831) );
  OAI21X1 U596 ( .A(n5571), .B(n3513), .C(n5832), .Y(n8588) );
  NAND2X1 U597 ( .A(arr[286]), .B(n3516), .Y(n5832) );
  NAND2X1 U598 ( .A(n5748), .B(n5660), .Y(n5791) );
  OAI21X1 U599 ( .A(n5491), .B(n3507), .C(n5834), .Y(n8589) );
  NAND2X1 U600 ( .A(arr[287]), .B(n3510), .Y(n5834) );
  OAI21X1 U601 ( .A(n5493), .B(n3507), .C(n5835), .Y(n8590) );
  NAND2X1 U602 ( .A(arr[288]), .B(n3510), .Y(n5835) );
  OAI21X1 U603 ( .A(n5495), .B(n3507), .C(n5836), .Y(n8591) );
  NAND2X1 U604 ( .A(arr[289]), .B(n3510), .Y(n5836) );
  OAI21X1 U605 ( .A(n5497), .B(n3507), .C(n5837), .Y(n8592) );
  NAND2X1 U606 ( .A(arr[290]), .B(n3510), .Y(n5837) );
  OAI21X1 U607 ( .A(n5499), .B(n3507), .C(n5838), .Y(n8593) );
  NAND2X1 U608 ( .A(arr[291]), .B(n3510), .Y(n5838) );
  OAI21X1 U609 ( .A(n5501), .B(n3508), .C(n5839), .Y(n8594) );
  NAND2X1 U610 ( .A(arr[292]), .B(n3510), .Y(n5839) );
  OAI21X1 U611 ( .A(n5503), .B(n3508), .C(n5840), .Y(n8595) );
  NAND2X1 U612 ( .A(arr[293]), .B(n3510), .Y(n5840) );
  OAI21X1 U613 ( .A(n5505), .B(n3508), .C(n5841), .Y(n8596) );
  NAND2X1 U614 ( .A(arr[294]), .B(n3510), .Y(n5841) );
  OAI21X1 U615 ( .A(n5507), .B(n3507), .C(n5842), .Y(n8597) );
  NAND2X1 U616 ( .A(arr[295]), .B(n3510), .Y(n5842) );
  OAI21X1 U617 ( .A(n5509), .B(n3508), .C(n5843), .Y(n8598) );
  NAND2X1 U618 ( .A(arr[296]), .B(n3510), .Y(n5843) );
  OAI21X1 U619 ( .A(n5511), .B(n3509), .C(n5844), .Y(n8599) );
  NAND2X1 U620 ( .A(arr[297]), .B(n3510), .Y(n5844) );
  OAI21X1 U621 ( .A(n5513), .B(n3509), .C(n5845), .Y(n8600) );
  NAND2X1 U622 ( .A(arr[298]), .B(n3510), .Y(n5845) );
  OAI21X1 U623 ( .A(n5515), .B(n3509), .C(n5846), .Y(n8601) );
  NAND2X1 U624 ( .A(arr[299]), .B(n3510), .Y(n5846) );
  OAI21X1 U625 ( .A(n5517), .B(n3508), .C(n5847), .Y(n8602) );
  NAND2X1 U626 ( .A(arr[300]), .B(n3511), .Y(n5847) );
  OAI21X1 U627 ( .A(n5519), .B(n3510), .C(n5848), .Y(n8603) );
  NAND2X1 U628 ( .A(arr[301]), .B(n3511), .Y(n5848) );
  OAI21X1 U629 ( .A(n5521), .B(n3510), .C(n5849), .Y(n8604) );
  NAND2X1 U630 ( .A(arr[302]), .B(n3511), .Y(n5849) );
  OAI21X1 U631 ( .A(n5523), .B(n3509), .C(n5850), .Y(n8605) );
  NAND2X1 U632 ( .A(arr[303]), .B(n3511), .Y(n5850) );
  OAI21X1 U633 ( .A(n5525), .B(n3509), .C(n5851), .Y(n8606) );
  NAND2X1 U634 ( .A(arr[304]), .B(n3511), .Y(n5851) );
  OAI21X1 U635 ( .A(n5527), .B(n3509), .C(n5852), .Y(n8607) );
  NAND2X1 U636 ( .A(arr[305]), .B(n3511), .Y(n5852) );
  OAI21X1 U637 ( .A(n5529), .B(n3509), .C(n5853), .Y(n8608) );
  NAND2X1 U638 ( .A(arr[306]), .B(n3511), .Y(n5853) );
  OAI21X1 U639 ( .A(n5531), .B(n3509), .C(n5854), .Y(n8609) );
  NAND2X1 U640 ( .A(arr[307]), .B(n3511), .Y(n5854) );
  OAI21X1 U641 ( .A(n5533), .B(n3509), .C(n5855), .Y(n8610) );
  NAND2X1 U642 ( .A(arr[308]), .B(n3511), .Y(n5855) );
  OAI21X1 U643 ( .A(n5535), .B(n3509), .C(n5856), .Y(n8611) );
  NAND2X1 U644 ( .A(arr[309]), .B(n3511), .Y(n5856) );
  OAI21X1 U645 ( .A(n5537), .B(n3509), .C(n5857), .Y(n8612) );
  NAND2X1 U646 ( .A(arr[310]), .B(n3511), .Y(n5857) );
  OAI21X1 U647 ( .A(n5539), .B(n3509), .C(n5858), .Y(n8613) );
  NAND2X1 U648 ( .A(arr[311]), .B(n3511), .Y(n5858) );
  OAI21X1 U649 ( .A(n5541), .B(n3509), .C(n5859), .Y(n8614) );
  NAND2X1 U650 ( .A(arr[312]), .B(n3511), .Y(n5859) );
  OAI21X1 U651 ( .A(n5543), .B(n3508), .C(n5860), .Y(n8615) );
  NAND2X1 U652 ( .A(arr[313]), .B(n3511), .Y(n5860) );
  OAI21X1 U653 ( .A(n5545), .B(n3508), .C(n5861), .Y(n8616) );
  NAND2X1 U654 ( .A(arr[314]), .B(n3511), .Y(n5861) );
  OAI21X1 U655 ( .A(n5547), .B(n3508), .C(n5862), .Y(n8617) );
  NAND2X1 U656 ( .A(arr[315]), .B(n3511), .Y(n5862) );
  OAI21X1 U657 ( .A(n5549), .B(n3508), .C(n5863), .Y(n8618) );
  NAND2X1 U658 ( .A(arr[316]), .B(n3511), .Y(n5863) );
  OAI21X1 U659 ( .A(n5551), .B(n3508), .C(n5864), .Y(n8619) );
  NAND2X1 U660 ( .A(arr[317]), .B(n3512), .Y(n5864) );
  OAI21X1 U661 ( .A(n5553), .B(n3508), .C(n5865), .Y(n8620) );
  NAND2X1 U662 ( .A(arr[318]), .B(n3512), .Y(n5865) );
  OAI21X1 U663 ( .A(n5555), .B(n3508), .C(n5866), .Y(n8621) );
  NAND2X1 U664 ( .A(arr[319]), .B(n3512), .Y(n5866) );
  OAI21X1 U665 ( .A(n5557), .B(n3508), .C(n5867), .Y(n8622) );
  NAND2X1 U666 ( .A(arr[320]), .B(n3512), .Y(n5867) );
  OAI21X1 U667 ( .A(n5559), .B(n3507), .C(n5868), .Y(n8623) );
  NAND2X1 U668 ( .A(arr[321]), .B(n3512), .Y(n5868) );
  OAI21X1 U669 ( .A(n5561), .B(n3507), .C(n5869), .Y(n8624) );
  NAND2X1 U670 ( .A(arr[322]), .B(n3512), .Y(n5869) );
  OAI21X1 U671 ( .A(n5563), .B(n3507), .C(n5870), .Y(n8625) );
  NAND2X1 U672 ( .A(arr[323]), .B(n3512), .Y(n5870) );
  OAI21X1 U673 ( .A(n5565), .B(n3507), .C(n5871), .Y(n8626) );
  NAND2X1 U674 ( .A(arr[324]), .B(n3512), .Y(n5871) );
  OAI21X1 U675 ( .A(n5567), .B(n3507), .C(n5872), .Y(n8627) );
  NAND2X1 U676 ( .A(arr[325]), .B(n3512), .Y(n5872) );
  OAI21X1 U677 ( .A(n5569), .B(n3507), .C(n5873), .Y(n8628) );
  NAND2X1 U678 ( .A(arr[326]), .B(n3510), .Y(n5873) );
  OAI21X1 U679 ( .A(n5571), .B(n3507), .C(n5874), .Y(n8629) );
  NAND2X1 U680 ( .A(arr[327]), .B(n3510), .Y(n5874) );
  NAND2X1 U681 ( .A(n5748), .B(n5703), .Y(n5833) );
  OAI21X1 U683 ( .A(n5491), .B(n3501), .C(n5877), .Y(n8630) );
  NAND2X1 U684 ( .A(arr[328]), .B(n3504), .Y(n5877) );
  OAI21X1 U685 ( .A(n5493), .B(n3501), .C(n5878), .Y(n8631) );
  NAND2X1 U686 ( .A(arr[329]), .B(n3504), .Y(n5878) );
  OAI21X1 U687 ( .A(n5495), .B(n3501), .C(n5879), .Y(n8632) );
  NAND2X1 U688 ( .A(arr[330]), .B(n3504), .Y(n5879) );
  OAI21X1 U689 ( .A(n5497), .B(n3501), .C(n5880), .Y(n8633) );
  NAND2X1 U690 ( .A(arr[331]), .B(n3504), .Y(n5880) );
  OAI21X1 U691 ( .A(n5499), .B(n3501), .C(n5881), .Y(n8634) );
  NAND2X1 U692 ( .A(arr[332]), .B(n3504), .Y(n5881) );
  OAI21X1 U693 ( .A(n5501), .B(n3502), .C(n5882), .Y(n8635) );
  NAND2X1 U694 ( .A(arr[333]), .B(n3504), .Y(n5882) );
  OAI21X1 U695 ( .A(n5503), .B(n3502), .C(n5883), .Y(n8636) );
  NAND2X1 U696 ( .A(arr[334]), .B(n3504), .Y(n5883) );
  OAI21X1 U697 ( .A(n5505), .B(n3502), .C(n5884), .Y(n8637) );
  NAND2X1 U698 ( .A(arr[335]), .B(n3504), .Y(n5884) );
  OAI21X1 U699 ( .A(n5507), .B(n3501), .C(n5885), .Y(n8638) );
  NAND2X1 U700 ( .A(arr[336]), .B(n3504), .Y(n5885) );
  OAI21X1 U701 ( .A(n5509), .B(n3502), .C(n5886), .Y(n8639) );
  NAND2X1 U702 ( .A(arr[337]), .B(n3504), .Y(n5886) );
  OAI21X1 U703 ( .A(n5511), .B(n3503), .C(n5887), .Y(n8640) );
  NAND2X1 U704 ( .A(arr[338]), .B(n3504), .Y(n5887) );
  OAI21X1 U705 ( .A(n5513), .B(n3503), .C(n5888), .Y(n8641) );
  NAND2X1 U706 ( .A(arr[339]), .B(n3504), .Y(n5888) );
  OAI21X1 U707 ( .A(n5515), .B(n3503), .C(n5889), .Y(n8642) );
  NAND2X1 U708 ( .A(arr[340]), .B(n3504), .Y(n5889) );
  OAI21X1 U709 ( .A(n5517), .B(n3502), .C(n5890), .Y(n8643) );
  NAND2X1 U710 ( .A(arr[341]), .B(n3505), .Y(n5890) );
  OAI21X1 U711 ( .A(n5519), .B(n3504), .C(n5891), .Y(n8644) );
  NAND2X1 U712 ( .A(arr[342]), .B(n3505), .Y(n5891) );
  OAI21X1 U713 ( .A(n5521), .B(n3504), .C(n5892), .Y(n8645) );
  NAND2X1 U714 ( .A(arr[343]), .B(n3505), .Y(n5892) );
  OAI21X1 U715 ( .A(n5523), .B(n3503), .C(n5893), .Y(n8646) );
  NAND2X1 U716 ( .A(arr[344]), .B(n3505), .Y(n5893) );
  OAI21X1 U717 ( .A(n5525), .B(n3503), .C(n5894), .Y(n8647) );
  NAND2X1 U718 ( .A(arr[345]), .B(n3505), .Y(n5894) );
  OAI21X1 U719 ( .A(n5527), .B(n3503), .C(n5895), .Y(n8648) );
  NAND2X1 U720 ( .A(arr[346]), .B(n3505), .Y(n5895) );
  OAI21X1 U721 ( .A(n5529), .B(n3503), .C(n5896), .Y(n8649) );
  NAND2X1 U722 ( .A(arr[347]), .B(n3505), .Y(n5896) );
  OAI21X1 U723 ( .A(n5531), .B(n3503), .C(n5897), .Y(n8650) );
  NAND2X1 U724 ( .A(arr[348]), .B(n3505), .Y(n5897) );
  OAI21X1 U725 ( .A(n5533), .B(n3503), .C(n5898), .Y(n8651) );
  NAND2X1 U726 ( .A(arr[349]), .B(n3505), .Y(n5898) );
  OAI21X1 U727 ( .A(n5535), .B(n3503), .C(n5899), .Y(n8652) );
  NAND2X1 U728 ( .A(arr[350]), .B(n3505), .Y(n5899) );
  OAI21X1 U729 ( .A(n5537), .B(n3503), .C(n5900), .Y(n8653) );
  NAND2X1 U730 ( .A(arr[351]), .B(n3505), .Y(n5900) );
  OAI21X1 U731 ( .A(n5539), .B(n3503), .C(n5901), .Y(n8654) );
  NAND2X1 U732 ( .A(arr[352]), .B(n3505), .Y(n5901) );
  OAI21X1 U733 ( .A(n5541), .B(n3503), .C(n5902), .Y(n8655) );
  NAND2X1 U734 ( .A(arr[353]), .B(n3505), .Y(n5902) );
  OAI21X1 U735 ( .A(n5543), .B(n3502), .C(n5903), .Y(n8656) );
  NAND2X1 U736 ( .A(arr[354]), .B(n3505), .Y(n5903) );
  OAI21X1 U737 ( .A(n5545), .B(n3502), .C(n5904), .Y(n8657) );
  NAND2X1 U738 ( .A(arr[355]), .B(n3505), .Y(n5904) );
  OAI21X1 U739 ( .A(n5547), .B(n3502), .C(n5905), .Y(n8658) );
  NAND2X1 U740 ( .A(arr[356]), .B(n3505), .Y(n5905) );
  OAI21X1 U741 ( .A(n5549), .B(n3502), .C(n5906), .Y(n8659) );
  NAND2X1 U742 ( .A(arr[357]), .B(n3505), .Y(n5906) );
  OAI21X1 U743 ( .A(n5551), .B(n3502), .C(n5907), .Y(n8660) );
  NAND2X1 U744 ( .A(arr[358]), .B(n3506), .Y(n5907) );
  OAI21X1 U745 ( .A(n5553), .B(n3502), .C(n5908), .Y(n8661) );
  NAND2X1 U746 ( .A(arr[359]), .B(n3506), .Y(n5908) );
  OAI21X1 U747 ( .A(n5555), .B(n3502), .C(n5909), .Y(n8662) );
  NAND2X1 U748 ( .A(arr[360]), .B(n3506), .Y(n5909) );
  OAI21X1 U749 ( .A(n5557), .B(n3502), .C(n5910), .Y(n8663) );
  NAND2X1 U750 ( .A(arr[361]), .B(n3506), .Y(n5910) );
  OAI21X1 U751 ( .A(n5559), .B(n3501), .C(n5911), .Y(n8664) );
  NAND2X1 U752 ( .A(arr[362]), .B(n3506), .Y(n5911) );
  OAI21X1 U753 ( .A(n5561), .B(n3501), .C(n5912), .Y(n8665) );
  NAND2X1 U754 ( .A(arr[363]), .B(n3506), .Y(n5912) );
  OAI21X1 U755 ( .A(n5563), .B(n3501), .C(n5913), .Y(n8666) );
  NAND2X1 U756 ( .A(arr[364]), .B(n3506), .Y(n5913) );
  OAI21X1 U757 ( .A(n5565), .B(n3501), .C(n5914), .Y(n8667) );
  NAND2X1 U758 ( .A(arr[365]), .B(n3506), .Y(n5914) );
  OAI21X1 U759 ( .A(n5567), .B(n3501), .C(n5915), .Y(n8668) );
  NAND2X1 U760 ( .A(arr[366]), .B(n3506), .Y(n5915) );
  OAI21X1 U761 ( .A(n5569), .B(n3501), .C(n5916), .Y(n8669) );
  NAND2X1 U762 ( .A(arr[367]), .B(n3504), .Y(n5916) );
  OAI21X1 U763 ( .A(n5571), .B(n3501), .C(n5917), .Y(n8670) );
  NAND2X1 U764 ( .A(arr[368]), .B(n3504), .Y(n5917) );
  NAND2X1 U765 ( .A(n5918), .B(n5573), .Y(n5876) );
  OAI21X1 U766 ( .A(n5491), .B(n3495), .C(n5920), .Y(n8671) );
  NAND2X1 U767 ( .A(arr[369]), .B(n3498), .Y(n5920) );
  OAI21X1 U768 ( .A(n5493), .B(n3495), .C(n5921), .Y(n8672) );
  NAND2X1 U769 ( .A(arr[370]), .B(n3498), .Y(n5921) );
  OAI21X1 U770 ( .A(n5495), .B(n3495), .C(n5922), .Y(n8673) );
  NAND2X1 U771 ( .A(arr[371]), .B(n3498), .Y(n5922) );
  OAI21X1 U772 ( .A(n5497), .B(n3495), .C(n5923), .Y(n8674) );
  NAND2X1 U773 ( .A(arr[372]), .B(n3498), .Y(n5923) );
  OAI21X1 U774 ( .A(n5499), .B(n3495), .C(n5924), .Y(n8675) );
  NAND2X1 U775 ( .A(arr[373]), .B(n3498), .Y(n5924) );
  OAI21X1 U776 ( .A(n5501), .B(n3496), .C(n5925), .Y(n8676) );
  NAND2X1 U777 ( .A(arr[374]), .B(n3498), .Y(n5925) );
  OAI21X1 U778 ( .A(n5503), .B(n3496), .C(n5926), .Y(n8677) );
  NAND2X1 U779 ( .A(arr[375]), .B(n3498), .Y(n5926) );
  OAI21X1 U780 ( .A(n5505), .B(n3496), .C(n5927), .Y(n8678) );
  NAND2X1 U781 ( .A(arr[376]), .B(n3498), .Y(n5927) );
  OAI21X1 U782 ( .A(n5507), .B(n3495), .C(n5928), .Y(n8679) );
  NAND2X1 U783 ( .A(arr[377]), .B(n3498), .Y(n5928) );
  OAI21X1 U784 ( .A(n5509), .B(n3496), .C(n5929), .Y(n8680) );
  NAND2X1 U785 ( .A(arr[378]), .B(n3498), .Y(n5929) );
  OAI21X1 U786 ( .A(n5511), .B(n3497), .C(n5930), .Y(n8681) );
  NAND2X1 U787 ( .A(arr[379]), .B(n3498), .Y(n5930) );
  OAI21X1 U788 ( .A(n5513), .B(n3497), .C(n5931), .Y(n8682) );
  NAND2X1 U789 ( .A(arr[380]), .B(n3498), .Y(n5931) );
  OAI21X1 U790 ( .A(n5515), .B(n3497), .C(n5932), .Y(n8683) );
  NAND2X1 U791 ( .A(arr[381]), .B(n3498), .Y(n5932) );
  OAI21X1 U792 ( .A(n5517), .B(n3496), .C(n5933), .Y(n8684) );
  NAND2X1 U793 ( .A(arr[382]), .B(n3499), .Y(n5933) );
  OAI21X1 U794 ( .A(n5519), .B(n3498), .C(n5934), .Y(n8685) );
  NAND2X1 U795 ( .A(arr[383]), .B(n3499), .Y(n5934) );
  OAI21X1 U796 ( .A(n5521), .B(n3498), .C(n5935), .Y(n8686) );
  NAND2X1 U797 ( .A(arr[384]), .B(n3499), .Y(n5935) );
  OAI21X1 U798 ( .A(n5523), .B(n3497), .C(n5936), .Y(n8687) );
  NAND2X1 U799 ( .A(arr[385]), .B(n3499), .Y(n5936) );
  OAI21X1 U800 ( .A(n5525), .B(n3497), .C(n5937), .Y(n8688) );
  NAND2X1 U801 ( .A(arr[386]), .B(n3499), .Y(n5937) );
  OAI21X1 U802 ( .A(n5527), .B(n3497), .C(n5938), .Y(n8689) );
  NAND2X1 U803 ( .A(arr[387]), .B(n3499), .Y(n5938) );
  OAI21X1 U804 ( .A(n5529), .B(n3497), .C(n5939), .Y(n8690) );
  NAND2X1 U805 ( .A(arr[388]), .B(n3499), .Y(n5939) );
  OAI21X1 U806 ( .A(n5531), .B(n3497), .C(n5940), .Y(n8691) );
  NAND2X1 U807 ( .A(arr[389]), .B(n3499), .Y(n5940) );
  OAI21X1 U808 ( .A(n5533), .B(n3497), .C(n5941), .Y(n8692) );
  NAND2X1 U809 ( .A(arr[390]), .B(n3499), .Y(n5941) );
  OAI21X1 U810 ( .A(n5535), .B(n3497), .C(n5942), .Y(n8693) );
  NAND2X1 U811 ( .A(arr[391]), .B(n3499), .Y(n5942) );
  OAI21X1 U812 ( .A(n5537), .B(n3497), .C(n5943), .Y(n8694) );
  NAND2X1 U813 ( .A(arr[392]), .B(n3499), .Y(n5943) );
  OAI21X1 U814 ( .A(n5539), .B(n3497), .C(n5944), .Y(n8695) );
  NAND2X1 U815 ( .A(arr[393]), .B(n3499), .Y(n5944) );
  OAI21X1 U816 ( .A(n5541), .B(n3497), .C(n5945), .Y(n8696) );
  NAND2X1 U817 ( .A(arr[394]), .B(n3499), .Y(n5945) );
  OAI21X1 U818 ( .A(n5543), .B(n3496), .C(n5946), .Y(n8697) );
  NAND2X1 U819 ( .A(arr[395]), .B(n3499), .Y(n5946) );
  OAI21X1 U820 ( .A(n5545), .B(n3496), .C(n5947), .Y(n8698) );
  NAND2X1 U821 ( .A(arr[396]), .B(n3499), .Y(n5947) );
  OAI21X1 U822 ( .A(n5547), .B(n3496), .C(n5948), .Y(n8699) );
  NAND2X1 U823 ( .A(arr[397]), .B(n3499), .Y(n5948) );
  OAI21X1 U824 ( .A(n5549), .B(n3496), .C(n5949), .Y(n8700) );
  NAND2X1 U825 ( .A(arr[398]), .B(n3499), .Y(n5949) );
  OAI21X1 U826 ( .A(n5551), .B(n3496), .C(n5950), .Y(n8701) );
  NAND2X1 U827 ( .A(arr[399]), .B(n3500), .Y(n5950) );
  OAI21X1 U828 ( .A(n5553), .B(n3496), .C(n5951), .Y(n8702) );
  NAND2X1 U829 ( .A(arr[400]), .B(n3500), .Y(n5951) );
  OAI21X1 U830 ( .A(n5555), .B(n3496), .C(n5952), .Y(n8703) );
  NAND2X1 U831 ( .A(arr[401]), .B(n3500), .Y(n5952) );
  OAI21X1 U832 ( .A(n5557), .B(n3496), .C(n5953), .Y(n8704) );
  NAND2X1 U833 ( .A(arr[402]), .B(n3500), .Y(n5953) );
  OAI21X1 U834 ( .A(n5559), .B(n3495), .C(n5954), .Y(n8705) );
  NAND2X1 U835 ( .A(arr[403]), .B(n3500), .Y(n5954) );
  OAI21X1 U836 ( .A(n5561), .B(n3495), .C(n5955), .Y(n8706) );
  NAND2X1 U837 ( .A(arr[404]), .B(n3500), .Y(n5955) );
  OAI21X1 U838 ( .A(n5563), .B(n3495), .C(n5956), .Y(n8707) );
  NAND2X1 U839 ( .A(arr[405]), .B(n3500), .Y(n5956) );
  OAI21X1 U840 ( .A(n5565), .B(n3495), .C(n5957), .Y(n8708) );
  NAND2X1 U841 ( .A(arr[406]), .B(n3500), .Y(n5957) );
  OAI21X1 U842 ( .A(n5567), .B(n3495), .C(n5958), .Y(n8709) );
  NAND2X1 U843 ( .A(arr[407]), .B(n3500), .Y(n5958) );
  OAI21X1 U844 ( .A(n5569), .B(n3495), .C(n5959), .Y(n8710) );
  NAND2X1 U845 ( .A(arr[408]), .B(n3498), .Y(n5959) );
  OAI21X1 U846 ( .A(n5571), .B(n3495), .C(n5960), .Y(n8711) );
  NAND2X1 U847 ( .A(arr[409]), .B(n3498), .Y(n5960) );
  NAND2X1 U848 ( .A(n5918), .B(n5617), .Y(n5919) );
  OAI21X1 U849 ( .A(n5491), .B(n3489), .C(n5962), .Y(n8712) );
  NAND2X1 U850 ( .A(arr[410]), .B(n3492), .Y(n5962) );
  OAI21X1 U851 ( .A(n5493), .B(n3489), .C(n5963), .Y(n8713) );
  NAND2X1 U852 ( .A(arr[411]), .B(n3492), .Y(n5963) );
  OAI21X1 U853 ( .A(n5495), .B(n3489), .C(n5964), .Y(n8714) );
  NAND2X1 U854 ( .A(arr[412]), .B(n3492), .Y(n5964) );
  OAI21X1 U855 ( .A(n5497), .B(n3489), .C(n5965), .Y(n8715) );
  NAND2X1 U856 ( .A(arr[413]), .B(n3492), .Y(n5965) );
  OAI21X1 U857 ( .A(n5499), .B(n3489), .C(n5966), .Y(n8716) );
  NAND2X1 U858 ( .A(arr[414]), .B(n3492), .Y(n5966) );
  OAI21X1 U859 ( .A(n5501), .B(n3490), .C(n5967), .Y(n8717) );
  NAND2X1 U860 ( .A(arr[415]), .B(n3492), .Y(n5967) );
  OAI21X1 U861 ( .A(n5503), .B(n3490), .C(n5968), .Y(n8718) );
  NAND2X1 U862 ( .A(arr[416]), .B(n3492), .Y(n5968) );
  OAI21X1 U863 ( .A(n5505), .B(n3490), .C(n5969), .Y(n8719) );
  NAND2X1 U864 ( .A(arr[417]), .B(n3492), .Y(n5969) );
  OAI21X1 U865 ( .A(n5507), .B(n3489), .C(n5970), .Y(n8720) );
  NAND2X1 U866 ( .A(arr[418]), .B(n3492), .Y(n5970) );
  OAI21X1 U867 ( .A(n5509), .B(n3490), .C(n5971), .Y(n8721) );
  NAND2X1 U868 ( .A(arr[419]), .B(n3492), .Y(n5971) );
  OAI21X1 U869 ( .A(n5511), .B(n3491), .C(n5972), .Y(n8722) );
  NAND2X1 U870 ( .A(arr[420]), .B(n3492), .Y(n5972) );
  OAI21X1 U871 ( .A(n5513), .B(n3491), .C(n5973), .Y(n8723) );
  NAND2X1 U872 ( .A(arr[421]), .B(n3492), .Y(n5973) );
  OAI21X1 U873 ( .A(n5515), .B(n3491), .C(n5974), .Y(n8724) );
  NAND2X1 U874 ( .A(arr[422]), .B(n3492), .Y(n5974) );
  OAI21X1 U875 ( .A(n5517), .B(n3490), .C(n5975), .Y(n8725) );
  NAND2X1 U876 ( .A(arr[423]), .B(n3493), .Y(n5975) );
  OAI21X1 U877 ( .A(n5519), .B(n3492), .C(n5976), .Y(n8726) );
  NAND2X1 U878 ( .A(arr[424]), .B(n3493), .Y(n5976) );
  OAI21X1 U879 ( .A(n5521), .B(n3492), .C(n5977), .Y(n8727) );
  NAND2X1 U880 ( .A(arr[425]), .B(n3493), .Y(n5977) );
  OAI21X1 U881 ( .A(n5523), .B(n3491), .C(n5978), .Y(n8728) );
  NAND2X1 U882 ( .A(arr[426]), .B(n3493), .Y(n5978) );
  OAI21X1 U883 ( .A(n5525), .B(n3491), .C(n5979), .Y(n8729) );
  NAND2X1 U884 ( .A(arr[427]), .B(n3493), .Y(n5979) );
  OAI21X1 U885 ( .A(n5527), .B(n3491), .C(n5980), .Y(n8730) );
  NAND2X1 U886 ( .A(arr[428]), .B(n3493), .Y(n5980) );
  OAI21X1 U887 ( .A(n5529), .B(n3491), .C(n5981), .Y(n8731) );
  NAND2X1 U888 ( .A(arr[429]), .B(n3493), .Y(n5981) );
  OAI21X1 U889 ( .A(n5531), .B(n3491), .C(n5982), .Y(n8732) );
  NAND2X1 U890 ( .A(arr[430]), .B(n3493), .Y(n5982) );
  OAI21X1 U891 ( .A(n5533), .B(n3491), .C(n5983), .Y(n8733) );
  NAND2X1 U892 ( .A(arr[431]), .B(n3493), .Y(n5983) );
  OAI21X1 U893 ( .A(n5535), .B(n3491), .C(n5984), .Y(n8734) );
  NAND2X1 U894 ( .A(arr[432]), .B(n3493), .Y(n5984) );
  OAI21X1 U895 ( .A(n5537), .B(n3491), .C(n5985), .Y(n8735) );
  NAND2X1 U896 ( .A(arr[433]), .B(n3493), .Y(n5985) );
  OAI21X1 U897 ( .A(n5539), .B(n3491), .C(n5986), .Y(n8736) );
  NAND2X1 U898 ( .A(arr[434]), .B(n3493), .Y(n5986) );
  OAI21X1 U899 ( .A(n5541), .B(n3491), .C(n5987), .Y(n8737) );
  NAND2X1 U900 ( .A(arr[435]), .B(n3493), .Y(n5987) );
  OAI21X1 U901 ( .A(n5543), .B(n3490), .C(n5988), .Y(n8738) );
  NAND2X1 U902 ( .A(arr[436]), .B(n3493), .Y(n5988) );
  OAI21X1 U903 ( .A(n5545), .B(n3490), .C(n5989), .Y(n8739) );
  NAND2X1 U904 ( .A(arr[437]), .B(n3493), .Y(n5989) );
  OAI21X1 U905 ( .A(n5547), .B(n3490), .C(n5990), .Y(n8740) );
  NAND2X1 U906 ( .A(arr[438]), .B(n3493), .Y(n5990) );
  OAI21X1 U907 ( .A(n5549), .B(n3490), .C(n5991), .Y(n8741) );
  NAND2X1 U908 ( .A(arr[439]), .B(n3493), .Y(n5991) );
  OAI21X1 U909 ( .A(n5551), .B(n3490), .C(n5992), .Y(n8742) );
  NAND2X1 U910 ( .A(arr[440]), .B(n3494), .Y(n5992) );
  OAI21X1 U911 ( .A(n5553), .B(n3490), .C(n5993), .Y(n8743) );
  NAND2X1 U912 ( .A(arr[441]), .B(n3494), .Y(n5993) );
  OAI21X1 U913 ( .A(n5555), .B(n3490), .C(n5994), .Y(n8744) );
  NAND2X1 U914 ( .A(arr[442]), .B(n3494), .Y(n5994) );
  OAI21X1 U915 ( .A(n5557), .B(n3490), .C(n5995), .Y(n8745) );
  NAND2X1 U916 ( .A(arr[443]), .B(n3494), .Y(n5995) );
  OAI21X1 U917 ( .A(n5559), .B(n3489), .C(n5996), .Y(n8746) );
  NAND2X1 U918 ( .A(arr[444]), .B(n3494), .Y(n5996) );
  OAI21X1 U919 ( .A(n5561), .B(n3489), .C(n5997), .Y(n8747) );
  NAND2X1 U920 ( .A(arr[445]), .B(n3494), .Y(n5997) );
  OAI21X1 U921 ( .A(n5563), .B(n3489), .C(n5998), .Y(n8748) );
  NAND2X1 U922 ( .A(arr[446]), .B(n3494), .Y(n5998) );
  OAI21X1 U923 ( .A(n5565), .B(n3489), .C(n5999), .Y(n8749) );
  NAND2X1 U924 ( .A(arr[447]), .B(n3494), .Y(n5999) );
  OAI21X1 U925 ( .A(n5567), .B(n3489), .C(n6000), .Y(n8750) );
  NAND2X1 U926 ( .A(arr[448]), .B(n3494), .Y(n6000) );
  OAI21X1 U927 ( .A(n5569), .B(n3489), .C(n6001), .Y(n8751) );
  NAND2X1 U928 ( .A(arr[449]), .B(n3492), .Y(n6001) );
  OAI21X1 U929 ( .A(n5571), .B(n3489), .C(n6002), .Y(n8752) );
  NAND2X1 U930 ( .A(arr[450]), .B(n3492), .Y(n6002) );
  NAND2X1 U931 ( .A(n5918), .B(n5660), .Y(n5961) );
  OAI21X1 U932 ( .A(n5491), .B(n3483), .C(n6004), .Y(n8753) );
  NAND2X1 U933 ( .A(arr[451]), .B(n3486), .Y(n6004) );
  OAI21X1 U934 ( .A(n5493), .B(n3483), .C(n6005), .Y(n8754) );
  NAND2X1 U935 ( .A(arr[452]), .B(n3486), .Y(n6005) );
  OAI21X1 U936 ( .A(n5495), .B(n3483), .C(n6006), .Y(n8755) );
  NAND2X1 U937 ( .A(arr[453]), .B(n3486), .Y(n6006) );
  OAI21X1 U938 ( .A(n5497), .B(n3483), .C(n6007), .Y(n8756) );
  NAND2X1 U939 ( .A(arr[454]), .B(n3486), .Y(n6007) );
  OAI21X1 U940 ( .A(n5499), .B(n3483), .C(n6008), .Y(n8757) );
  NAND2X1 U941 ( .A(arr[455]), .B(n3486), .Y(n6008) );
  OAI21X1 U942 ( .A(n5501), .B(n3484), .C(n6009), .Y(n8758) );
  NAND2X1 U943 ( .A(arr[456]), .B(n3486), .Y(n6009) );
  OAI21X1 U944 ( .A(n5503), .B(n3484), .C(n6010), .Y(n8759) );
  NAND2X1 U945 ( .A(arr[457]), .B(n3486), .Y(n6010) );
  OAI21X1 U946 ( .A(n5505), .B(n3484), .C(n6011), .Y(n8760) );
  NAND2X1 U947 ( .A(arr[458]), .B(n3486), .Y(n6011) );
  OAI21X1 U948 ( .A(n5507), .B(n3483), .C(n6012), .Y(n8761) );
  NAND2X1 U949 ( .A(arr[459]), .B(n3486), .Y(n6012) );
  OAI21X1 U950 ( .A(n5509), .B(n3484), .C(n6013), .Y(n8762) );
  NAND2X1 U951 ( .A(arr[460]), .B(n3486), .Y(n6013) );
  OAI21X1 U952 ( .A(n5511), .B(n3485), .C(n6014), .Y(n8763) );
  NAND2X1 U953 ( .A(arr[461]), .B(n3486), .Y(n6014) );
  OAI21X1 U954 ( .A(n5513), .B(n3485), .C(n6015), .Y(n8764) );
  NAND2X1 U955 ( .A(arr[462]), .B(n3486), .Y(n6015) );
  OAI21X1 U956 ( .A(n5515), .B(n3485), .C(n6016), .Y(n8765) );
  NAND2X1 U957 ( .A(arr[463]), .B(n3486), .Y(n6016) );
  OAI21X1 U958 ( .A(n5517), .B(n3484), .C(n6017), .Y(n8766) );
  NAND2X1 U959 ( .A(arr[464]), .B(n3487), .Y(n6017) );
  OAI21X1 U960 ( .A(n5519), .B(n3486), .C(n6018), .Y(n8767) );
  NAND2X1 U961 ( .A(arr[465]), .B(n3487), .Y(n6018) );
  OAI21X1 U962 ( .A(n5521), .B(n3486), .C(n6019), .Y(n8768) );
  NAND2X1 U963 ( .A(arr[466]), .B(n3487), .Y(n6019) );
  OAI21X1 U964 ( .A(n5523), .B(n3485), .C(n6020), .Y(n8769) );
  NAND2X1 U965 ( .A(arr[467]), .B(n3487), .Y(n6020) );
  OAI21X1 U966 ( .A(n5525), .B(n3485), .C(n6021), .Y(n8770) );
  NAND2X1 U967 ( .A(arr[468]), .B(n3487), .Y(n6021) );
  OAI21X1 U968 ( .A(n5527), .B(n3485), .C(n6022), .Y(n8771) );
  NAND2X1 U969 ( .A(arr[469]), .B(n3487), .Y(n6022) );
  OAI21X1 U970 ( .A(n5529), .B(n3485), .C(n6023), .Y(n8772) );
  NAND2X1 U971 ( .A(arr[470]), .B(n3487), .Y(n6023) );
  OAI21X1 U972 ( .A(n5531), .B(n3485), .C(n6024), .Y(n8773) );
  NAND2X1 U973 ( .A(arr[471]), .B(n3487), .Y(n6024) );
  OAI21X1 U974 ( .A(n5533), .B(n3485), .C(n6025), .Y(n8774) );
  NAND2X1 U975 ( .A(arr[472]), .B(n3487), .Y(n6025) );
  OAI21X1 U976 ( .A(n5535), .B(n3485), .C(n6026), .Y(n8775) );
  NAND2X1 U977 ( .A(arr[473]), .B(n3487), .Y(n6026) );
  OAI21X1 U978 ( .A(n5537), .B(n3485), .C(n6027), .Y(n8776) );
  NAND2X1 U979 ( .A(arr[474]), .B(n3487), .Y(n6027) );
  OAI21X1 U980 ( .A(n5539), .B(n3485), .C(n6028), .Y(n8777) );
  NAND2X1 U981 ( .A(arr[475]), .B(n3487), .Y(n6028) );
  OAI21X1 U982 ( .A(n5541), .B(n3485), .C(n6029), .Y(n8778) );
  NAND2X1 U983 ( .A(arr[476]), .B(n3487), .Y(n6029) );
  OAI21X1 U984 ( .A(n5543), .B(n3484), .C(n6030), .Y(n8779) );
  NAND2X1 U985 ( .A(arr[477]), .B(n3487), .Y(n6030) );
  OAI21X1 U986 ( .A(n5545), .B(n3484), .C(n6031), .Y(n8780) );
  NAND2X1 U987 ( .A(arr[478]), .B(n3487), .Y(n6031) );
  OAI21X1 U988 ( .A(n5547), .B(n3484), .C(n6032), .Y(n8781) );
  NAND2X1 U989 ( .A(arr[479]), .B(n3487), .Y(n6032) );
  OAI21X1 U990 ( .A(n5549), .B(n3484), .C(n6033), .Y(n8782) );
  NAND2X1 U991 ( .A(arr[480]), .B(n3487), .Y(n6033) );
  OAI21X1 U992 ( .A(n5551), .B(n3484), .C(n6034), .Y(n8783) );
  NAND2X1 U993 ( .A(arr[481]), .B(n3488), .Y(n6034) );
  OAI21X1 U994 ( .A(n5553), .B(n3484), .C(n6035), .Y(n8784) );
  NAND2X1 U995 ( .A(arr[482]), .B(n3488), .Y(n6035) );
  OAI21X1 U996 ( .A(n5555), .B(n3484), .C(n6036), .Y(n8785) );
  NAND2X1 U997 ( .A(arr[483]), .B(n3488), .Y(n6036) );
  OAI21X1 U998 ( .A(n5557), .B(n3484), .C(n6037), .Y(n8786) );
  NAND2X1 U999 ( .A(arr[484]), .B(n3488), .Y(n6037) );
  OAI21X1 U1000 ( .A(n5559), .B(n3483), .C(n6038), .Y(n8787) );
  NAND2X1 U1001 ( .A(arr[485]), .B(n3488), .Y(n6038) );
  OAI21X1 U1002 ( .A(n5561), .B(n3483), .C(n6039), .Y(n8788) );
  NAND2X1 U1003 ( .A(arr[486]), .B(n3488), .Y(n6039) );
  OAI21X1 U1004 ( .A(n5563), .B(n3483), .C(n6040), .Y(n8789) );
  NAND2X1 U1005 ( .A(arr[487]), .B(n3488), .Y(n6040) );
  OAI21X1 U1006 ( .A(n5565), .B(n3483), .C(n6041), .Y(n8790) );
  NAND2X1 U1007 ( .A(arr[488]), .B(n3488), .Y(n6041) );
  OAI21X1 U1008 ( .A(n5567), .B(n3483), .C(n6042), .Y(n8791) );
  NAND2X1 U1009 ( .A(arr[489]), .B(n3488), .Y(n6042) );
  OAI21X1 U1010 ( .A(n5569), .B(n3483), .C(n6043), .Y(n8792) );
  NAND2X1 U1011 ( .A(arr[490]), .B(n3486), .Y(n6043) );
  OAI21X1 U1012 ( .A(n5571), .B(n3483), .C(n6044), .Y(n8793) );
  NAND2X1 U1013 ( .A(arr[491]), .B(n3486), .Y(n6044) );
  NAND2X1 U1014 ( .A(n5918), .B(n5703), .Y(n6003) );
  OAI21X1 U1016 ( .A(n5491), .B(n3477), .C(n6047), .Y(n8794) );
  NAND2X1 U1017 ( .A(arr[492]), .B(n3480), .Y(n6047) );
  OAI21X1 U1018 ( .A(n5493), .B(n3477), .C(n6048), .Y(n8795) );
  NAND2X1 U1019 ( .A(arr[493]), .B(n3480), .Y(n6048) );
  OAI21X1 U1020 ( .A(n5495), .B(n3477), .C(n6049), .Y(n8796) );
  NAND2X1 U1021 ( .A(arr[494]), .B(n3480), .Y(n6049) );
  OAI21X1 U1022 ( .A(n5497), .B(n3477), .C(n6050), .Y(n8797) );
  NAND2X1 U1023 ( .A(arr[495]), .B(n3480), .Y(n6050) );
  OAI21X1 U1024 ( .A(n5499), .B(n3477), .C(n6051), .Y(n8798) );
  NAND2X1 U1025 ( .A(arr[496]), .B(n3480), .Y(n6051) );
  OAI21X1 U1026 ( .A(n5501), .B(n3478), .C(n6052), .Y(n8799) );
  NAND2X1 U1027 ( .A(arr[497]), .B(n3480), .Y(n6052) );
  OAI21X1 U1028 ( .A(n5503), .B(n3478), .C(n6053), .Y(n8800) );
  NAND2X1 U1029 ( .A(arr[498]), .B(n3480), .Y(n6053) );
  OAI21X1 U1030 ( .A(n5505), .B(n3478), .C(n6054), .Y(n8801) );
  NAND2X1 U1031 ( .A(arr[499]), .B(n3480), .Y(n6054) );
  OAI21X1 U1032 ( .A(n5507), .B(n3477), .C(n6055), .Y(n8802) );
  NAND2X1 U1033 ( .A(arr[500]), .B(n3480), .Y(n6055) );
  OAI21X1 U1034 ( .A(n5509), .B(n3478), .C(n6056), .Y(n8803) );
  NAND2X1 U1035 ( .A(arr[501]), .B(n3480), .Y(n6056) );
  OAI21X1 U1036 ( .A(n5511), .B(n3479), .C(n6057), .Y(n8804) );
  NAND2X1 U1037 ( .A(arr[502]), .B(n3480), .Y(n6057) );
  OAI21X1 U1038 ( .A(n5513), .B(n3479), .C(n6058), .Y(n8805) );
  NAND2X1 U1039 ( .A(arr[503]), .B(n3480), .Y(n6058) );
  OAI21X1 U1040 ( .A(n5515), .B(n3479), .C(n6059), .Y(n8806) );
  NAND2X1 U1041 ( .A(arr[504]), .B(n3480), .Y(n6059) );
  OAI21X1 U1042 ( .A(n5517), .B(n3478), .C(n6060), .Y(n8807) );
  NAND2X1 U1043 ( .A(arr[505]), .B(n3481), .Y(n6060) );
  OAI21X1 U1044 ( .A(n5519), .B(n3480), .C(n6061), .Y(n8808) );
  NAND2X1 U1045 ( .A(arr[506]), .B(n3481), .Y(n6061) );
  OAI21X1 U1046 ( .A(n5521), .B(n3480), .C(n6062), .Y(n8809) );
  NAND2X1 U1047 ( .A(arr[507]), .B(n3481), .Y(n6062) );
  OAI21X1 U1048 ( .A(n5523), .B(n3479), .C(n6063), .Y(n8810) );
  NAND2X1 U1049 ( .A(arr[508]), .B(n3481), .Y(n6063) );
  OAI21X1 U1050 ( .A(n5525), .B(n3479), .C(n6064), .Y(n8811) );
  NAND2X1 U1051 ( .A(arr[509]), .B(n3481), .Y(n6064) );
  OAI21X1 U1052 ( .A(n5527), .B(n3479), .C(n6065), .Y(n8812) );
  NAND2X1 U1053 ( .A(arr[510]), .B(n3481), .Y(n6065) );
  OAI21X1 U1054 ( .A(n5529), .B(n3479), .C(n6066), .Y(n8813) );
  NAND2X1 U1055 ( .A(arr[511]), .B(n3481), .Y(n6066) );
  OAI21X1 U1056 ( .A(n5531), .B(n3479), .C(n6067), .Y(n8814) );
  NAND2X1 U1057 ( .A(arr[512]), .B(n3481), .Y(n6067) );
  OAI21X1 U1058 ( .A(n5533), .B(n3479), .C(n6068), .Y(n8815) );
  NAND2X1 U1059 ( .A(arr[513]), .B(n3481), .Y(n6068) );
  OAI21X1 U1060 ( .A(n5535), .B(n3479), .C(n6069), .Y(n8816) );
  NAND2X1 U1061 ( .A(arr[514]), .B(n3481), .Y(n6069) );
  OAI21X1 U1062 ( .A(n5537), .B(n3479), .C(n6070), .Y(n8817) );
  NAND2X1 U1063 ( .A(arr[515]), .B(n3481), .Y(n6070) );
  OAI21X1 U1064 ( .A(n5539), .B(n3479), .C(n6071), .Y(n8818) );
  NAND2X1 U1065 ( .A(arr[516]), .B(n3481), .Y(n6071) );
  OAI21X1 U1066 ( .A(n5541), .B(n3479), .C(n6072), .Y(n8819) );
  NAND2X1 U1067 ( .A(arr[517]), .B(n3481), .Y(n6072) );
  OAI21X1 U1068 ( .A(n5543), .B(n3478), .C(n6073), .Y(n8820) );
  NAND2X1 U1069 ( .A(arr[518]), .B(n3481), .Y(n6073) );
  OAI21X1 U1070 ( .A(n5545), .B(n3478), .C(n6074), .Y(n8821) );
  NAND2X1 U1071 ( .A(arr[519]), .B(n3481), .Y(n6074) );
  OAI21X1 U1072 ( .A(n5547), .B(n3478), .C(n6075), .Y(n8822) );
  NAND2X1 U1073 ( .A(arr[520]), .B(n3481), .Y(n6075) );
  OAI21X1 U1074 ( .A(n5549), .B(n3478), .C(n6076), .Y(n8823) );
  NAND2X1 U1075 ( .A(arr[521]), .B(n3481), .Y(n6076) );
  OAI21X1 U1076 ( .A(n5551), .B(n3478), .C(n6077), .Y(n8824) );
  NAND2X1 U1077 ( .A(arr[522]), .B(n3482), .Y(n6077) );
  OAI21X1 U1078 ( .A(n5553), .B(n3478), .C(n6078), .Y(n8825) );
  NAND2X1 U1079 ( .A(arr[523]), .B(n3482), .Y(n6078) );
  OAI21X1 U1080 ( .A(n5555), .B(n3478), .C(n6079), .Y(n8826) );
  NAND2X1 U1081 ( .A(arr[524]), .B(n3482), .Y(n6079) );
  OAI21X1 U1082 ( .A(n5557), .B(n3478), .C(n6080), .Y(n8827) );
  NAND2X1 U1083 ( .A(arr[525]), .B(n3482), .Y(n6080) );
  OAI21X1 U1084 ( .A(n5559), .B(n3477), .C(n6081), .Y(n8828) );
  NAND2X1 U1085 ( .A(arr[526]), .B(n3482), .Y(n6081) );
  OAI21X1 U1086 ( .A(n5561), .B(n3477), .C(n6082), .Y(n8829) );
  NAND2X1 U1087 ( .A(arr[527]), .B(n3482), .Y(n6082) );
  OAI21X1 U1088 ( .A(n5563), .B(n3477), .C(n6083), .Y(n8830) );
  NAND2X1 U1089 ( .A(arr[528]), .B(n3482), .Y(n6083) );
  OAI21X1 U1090 ( .A(n5565), .B(n3477), .C(n6084), .Y(n8831) );
  NAND2X1 U1091 ( .A(arr[529]), .B(n3482), .Y(n6084) );
  OAI21X1 U1092 ( .A(n5567), .B(n3477), .C(n6085), .Y(n8832) );
  NAND2X1 U1093 ( .A(arr[530]), .B(n3482), .Y(n6085) );
  OAI21X1 U1094 ( .A(n5569), .B(n3477), .C(n6086), .Y(n8833) );
  NAND2X1 U1095 ( .A(arr[531]), .B(n3480), .Y(n6086) );
  OAI21X1 U1096 ( .A(n5571), .B(n3477), .C(n6087), .Y(n8834) );
  NAND2X1 U1097 ( .A(arr[532]), .B(n3480), .Y(n6087) );
  NAND2X1 U1098 ( .A(n6088), .B(n5573), .Y(n6046) );
  OAI21X1 U1099 ( .A(n5491), .B(n3471), .C(n6090), .Y(n8835) );
  NAND2X1 U1100 ( .A(arr[533]), .B(n3474), .Y(n6090) );
  OAI21X1 U1101 ( .A(n5493), .B(n3471), .C(n6091), .Y(n8836) );
  NAND2X1 U1102 ( .A(arr[534]), .B(n3474), .Y(n6091) );
  OAI21X1 U1103 ( .A(n5495), .B(n3471), .C(n6092), .Y(n8837) );
  NAND2X1 U1104 ( .A(arr[535]), .B(n3474), .Y(n6092) );
  OAI21X1 U1105 ( .A(n5497), .B(n3471), .C(n6093), .Y(n8838) );
  NAND2X1 U1106 ( .A(arr[536]), .B(n3474), .Y(n6093) );
  OAI21X1 U1107 ( .A(n5499), .B(n3471), .C(n6094), .Y(n8839) );
  NAND2X1 U1108 ( .A(arr[537]), .B(n3474), .Y(n6094) );
  OAI21X1 U1109 ( .A(n5501), .B(n3472), .C(n6095), .Y(n8840) );
  NAND2X1 U1110 ( .A(arr[538]), .B(n3474), .Y(n6095) );
  OAI21X1 U1111 ( .A(n5503), .B(n3472), .C(n6096), .Y(n8841) );
  NAND2X1 U1112 ( .A(arr[539]), .B(n3474), .Y(n6096) );
  OAI21X1 U1113 ( .A(n5505), .B(n3472), .C(n6097), .Y(n8842) );
  NAND2X1 U1114 ( .A(arr[540]), .B(n3474), .Y(n6097) );
  OAI21X1 U1115 ( .A(n5507), .B(n3471), .C(n6098), .Y(n8843) );
  NAND2X1 U1116 ( .A(arr[541]), .B(n3474), .Y(n6098) );
  OAI21X1 U1117 ( .A(n5509), .B(n3472), .C(n6099), .Y(n8844) );
  NAND2X1 U1118 ( .A(arr[542]), .B(n3474), .Y(n6099) );
  OAI21X1 U1119 ( .A(n5511), .B(n3473), .C(n6100), .Y(n8845) );
  NAND2X1 U1120 ( .A(arr[543]), .B(n3474), .Y(n6100) );
  OAI21X1 U1121 ( .A(n5513), .B(n3473), .C(n6101), .Y(n8846) );
  NAND2X1 U1122 ( .A(arr[544]), .B(n3474), .Y(n6101) );
  OAI21X1 U1123 ( .A(n5515), .B(n3473), .C(n6102), .Y(n8847) );
  NAND2X1 U1124 ( .A(arr[545]), .B(n3474), .Y(n6102) );
  OAI21X1 U1125 ( .A(n5517), .B(n3472), .C(n6103), .Y(n8848) );
  NAND2X1 U1126 ( .A(arr[546]), .B(n3475), .Y(n6103) );
  OAI21X1 U1127 ( .A(n5519), .B(n3474), .C(n6104), .Y(n8849) );
  NAND2X1 U1128 ( .A(arr[547]), .B(n3475), .Y(n6104) );
  OAI21X1 U1129 ( .A(n5521), .B(n3474), .C(n6105), .Y(n8850) );
  NAND2X1 U1130 ( .A(arr[548]), .B(n3475), .Y(n6105) );
  OAI21X1 U1131 ( .A(n5523), .B(n3473), .C(n6106), .Y(n8851) );
  NAND2X1 U1132 ( .A(arr[549]), .B(n3475), .Y(n6106) );
  OAI21X1 U1133 ( .A(n5525), .B(n3473), .C(n6107), .Y(n8852) );
  NAND2X1 U1134 ( .A(arr[550]), .B(n3475), .Y(n6107) );
  OAI21X1 U1135 ( .A(n5527), .B(n3473), .C(n6108), .Y(n8853) );
  NAND2X1 U1136 ( .A(arr[551]), .B(n3475), .Y(n6108) );
  OAI21X1 U1137 ( .A(n5529), .B(n3473), .C(n6109), .Y(n8854) );
  NAND2X1 U1138 ( .A(arr[552]), .B(n3475), .Y(n6109) );
  OAI21X1 U1139 ( .A(n5531), .B(n3473), .C(n6110), .Y(n8855) );
  NAND2X1 U1140 ( .A(arr[553]), .B(n3475), .Y(n6110) );
  OAI21X1 U1141 ( .A(n5533), .B(n3473), .C(n6111), .Y(n8856) );
  NAND2X1 U1142 ( .A(arr[554]), .B(n3475), .Y(n6111) );
  OAI21X1 U1143 ( .A(n5535), .B(n3473), .C(n6112), .Y(n8857) );
  NAND2X1 U1144 ( .A(arr[555]), .B(n3475), .Y(n6112) );
  OAI21X1 U1145 ( .A(n5537), .B(n3473), .C(n6113), .Y(n8858) );
  NAND2X1 U1146 ( .A(arr[556]), .B(n3475), .Y(n6113) );
  OAI21X1 U1147 ( .A(n5539), .B(n3473), .C(n6114), .Y(n8859) );
  NAND2X1 U1148 ( .A(arr[557]), .B(n3475), .Y(n6114) );
  OAI21X1 U1149 ( .A(n5541), .B(n3473), .C(n6115), .Y(n8860) );
  NAND2X1 U1150 ( .A(arr[558]), .B(n3475), .Y(n6115) );
  OAI21X1 U1151 ( .A(n5543), .B(n3472), .C(n6116), .Y(n8861) );
  NAND2X1 U1152 ( .A(arr[559]), .B(n3475), .Y(n6116) );
  OAI21X1 U1153 ( .A(n5545), .B(n3472), .C(n6117), .Y(n8862) );
  NAND2X1 U1154 ( .A(arr[560]), .B(n3475), .Y(n6117) );
  OAI21X1 U1155 ( .A(n5547), .B(n3472), .C(n6118), .Y(n8863) );
  NAND2X1 U1156 ( .A(arr[561]), .B(n3475), .Y(n6118) );
  OAI21X1 U1157 ( .A(n5549), .B(n3472), .C(n6119), .Y(n8864) );
  NAND2X1 U1158 ( .A(arr[562]), .B(n3475), .Y(n6119) );
  OAI21X1 U1159 ( .A(n5551), .B(n3472), .C(n6120), .Y(n8865) );
  NAND2X1 U1160 ( .A(arr[563]), .B(n3476), .Y(n6120) );
  OAI21X1 U1161 ( .A(n5553), .B(n3472), .C(n6121), .Y(n8866) );
  NAND2X1 U1162 ( .A(arr[564]), .B(n3476), .Y(n6121) );
  OAI21X1 U1163 ( .A(n5555), .B(n3472), .C(n6122), .Y(n8867) );
  NAND2X1 U1164 ( .A(arr[565]), .B(n3476), .Y(n6122) );
  OAI21X1 U1165 ( .A(n5557), .B(n3472), .C(n6123), .Y(n8868) );
  NAND2X1 U1166 ( .A(arr[566]), .B(n3476), .Y(n6123) );
  OAI21X1 U1167 ( .A(n5559), .B(n3471), .C(n6124), .Y(n8869) );
  NAND2X1 U1168 ( .A(arr[567]), .B(n3476), .Y(n6124) );
  OAI21X1 U1169 ( .A(n5561), .B(n3471), .C(n6125), .Y(n8870) );
  NAND2X1 U1170 ( .A(arr[568]), .B(n3476), .Y(n6125) );
  OAI21X1 U1171 ( .A(n5563), .B(n3471), .C(n6126), .Y(n8871) );
  NAND2X1 U1172 ( .A(arr[569]), .B(n3476), .Y(n6126) );
  OAI21X1 U1173 ( .A(n5565), .B(n3471), .C(n6127), .Y(n8872) );
  NAND2X1 U1174 ( .A(arr[570]), .B(n3476), .Y(n6127) );
  OAI21X1 U1175 ( .A(n5567), .B(n3471), .C(n6128), .Y(n8873) );
  NAND2X1 U1176 ( .A(arr[571]), .B(n3476), .Y(n6128) );
  OAI21X1 U1177 ( .A(n5569), .B(n3471), .C(n6129), .Y(n8874) );
  NAND2X1 U1178 ( .A(arr[572]), .B(n3474), .Y(n6129) );
  OAI21X1 U1179 ( .A(n5571), .B(n3471), .C(n6130), .Y(n8875) );
  NAND2X1 U1180 ( .A(arr[573]), .B(n3474), .Y(n6130) );
  NAND2X1 U1181 ( .A(n6088), .B(n5617), .Y(n6089) );
  OAI21X1 U1182 ( .A(n5491), .B(n3465), .C(n6132), .Y(n8876) );
  NAND2X1 U1183 ( .A(arr[574]), .B(n3468), .Y(n6132) );
  OAI21X1 U1184 ( .A(n5493), .B(n3465), .C(n6133), .Y(n8877) );
  NAND2X1 U1185 ( .A(arr[575]), .B(n3468), .Y(n6133) );
  OAI21X1 U1186 ( .A(n5495), .B(n3465), .C(n6134), .Y(n8878) );
  NAND2X1 U1187 ( .A(arr[576]), .B(n3468), .Y(n6134) );
  OAI21X1 U1188 ( .A(n5497), .B(n3465), .C(n6135), .Y(n8879) );
  NAND2X1 U1189 ( .A(arr[577]), .B(n3468), .Y(n6135) );
  OAI21X1 U1190 ( .A(n5499), .B(n3465), .C(n6136), .Y(n8880) );
  NAND2X1 U1191 ( .A(arr[578]), .B(n3468), .Y(n6136) );
  OAI21X1 U1192 ( .A(n5501), .B(n3466), .C(n6137), .Y(n8881) );
  NAND2X1 U1193 ( .A(arr[579]), .B(n3468), .Y(n6137) );
  OAI21X1 U1194 ( .A(n5503), .B(n3466), .C(n6138), .Y(n8882) );
  NAND2X1 U1195 ( .A(arr[580]), .B(n3468), .Y(n6138) );
  OAI21X1 U1196 ( .A(n5505), .B(n3466), .C(n6139), .Y(n8883) );
  NAND2X1 U1197 ( .A(arr[581]), .B(n3468), .Y(n6139) );
  OAI21X1 U1198 ( .A(n5507), .B(n3465), .C(n6140), .Y(n8884) );
  NAND2X1 U1199 ( .A(arr[582]), .B(n3468), .Y(n6140) );
  OAI21X1 U1200 ( .A(n5509), .B(n3466), .C(n6141), .Y(n8885) );
  NAND2X1 U1201 ( .A(arr[583]), .B(n3468), .Y(n6141) );
  OAI21X1 U1202 ( .A(n5511), .B(n3467), .C(n6142), .Y(n8886) );
  NAND2X1 U1203 ( .A(arr[584]), .B(n3468), .Y(n6142) );
  OAI21X1 U1204 ( .A(n5513), .B(n3467), .C(n6143), .Y(n8887) );
  NAND2X1 U1205 ( .A(arr[585]), .B(n3468), .Y(n6143) );
  OAI21X1 U1206 ( .A(n5515), .B(n3467), .C(n6144), .Y(n8888) );
  NAND2X1 U1207 ( .A(arr[586]), .B(n3468), .Y(n6144) );
  OAI21X1 U1208 ( .A(n5517), .B(n3466), .C(n6145), .Y(n8889) );
  NAND2X1 U1209 ( .A(arr[587]), .B(n3469), .Y(n6145) );
  OAI21X1 U1210 ( .A(n5519), .B(n3468), .C(n6146), .Y(n8890) );
  NAND2X1 U1211 ( .A(arr[588]), .B(n3469), .Y(n6146) );
  OAI21X1 U1212 ( .A(n5521), .B(n3468), .C(n6147), .Y(n8891) );
  NAND2X1 U1213 ( .A(arr[589]), .B(n3469), .Y(n6147) );
  OAI21X1 U1214 ( .A(n5523), .B(n3467), .C(n6148), .Y(n8892) );
  NAND2X1 U1215 ( .A(arr[590]), .B(n3469), .Y(n6148) );
  OAI21X1 U1216 ( .A(n5525), .B(n3467), .C(n6149), .Y(n8893) );
  NAND2X1 U1217 ( .A(arr[591]), .B(n3469), .Y(n6149) );
  OAI21X1 U1218 ( .A(n5527), .B(n3467), .C(n6150), .Y(n8894) );
  NAND2X1 U1219 ( .A(arr[592]), .B(n3469), .Y(n6150) );
  OAI21X1 U1220 ( .A(n5529), .B(n3467), .C(n6151), .Y(n8895) );
  NAND2X1 U1221 ( .A(arr[593]), .B(n3469), .Y(n6151) );
  OAI21X1 U1222 ( .A(n5531), .B(n3467), .C(n6152), .Y(n8896) );
  NAND2X1 U1223 ( .A(arr[594]), .B(n3469), .Y(n6152) );
  OAI21X1 U1224 ( .A(n5533), .B(n3467), .C(n6153), .Y(n8897) );
  NAND2X1 U1225 ( .A(arr[595]), .B(n3469), .Y(n6153) );
  OAI21X1 U1226 ( .A(n5535), .B(n3467), .C(n6154), .Y(n8898) );
  NAND2X1 U1227 ( .A(arr[596]), .B(n3469), .Y(n6154) );
  OAI21X1 U1228 ( .A(n5537), .B(n3467), .C(n6155), .Y(n8899) );
  NAND2X1 U1229 ( .A(arr[597]), .B(n3469), .Y(n6155) );
  OAI21X1 U1230 ( .A(n5539), .B(n3467), .C(n6156), .Y(n8900) );
  NAND2X1 U1231 ( .A(arr[598]), .B(n3469), .Y(n6156) );
  OAI21X1 U1232 ( .A(n5541), .B(n3467), .C(n6157), .Y(n8901) );
  NAND2X1 U1233 ( .A(arr[599]), .B(n3469), .Y(n6157) );
  OAI21X1 U1234 ( .A(n5543), .B(n3466), .C(n6158), .Y(n8902) );
  NAND2X1 U1235 ( .A(arr[600]), .B(n3469), .Y(n6158) );
  OAI21X1 U1236 ( .A(n5545), .B(n3466), .C(n6159), .Y(n8903) );
  NAND2X1 U1237 ( .A(arr[601]), .B(n3469), .Y(n6159) );
  OAI21X1 U1238 ( .A(n5547), .B(n3466), .C(n6160), .Y(n8904) );
  NAND2X1 U1239 ( .A(arr[602]), .B(n3469), .Y(n6160) );
  OAI21X1 U1240 ( .A(n5549), .B(n3466), .C(n6161), .Y(n8905) );
  NAND2X1 U1241 ( .A(arr[603]), .B(n3469), .Y(n6161) );
  OAI21X1 U1242 ( .A(n5551), .B(n3466), .C(n6162), .Y(n8906) );
  NAND2X1 U1243 ( .A(arr[604]), .B(n3470), .Y(n6162) );
  OAI21X1 U1244 ( .A(n5553), .B(n3466), .C(n6163), .Y(n8907) );
  NAND2X1 U1245 ( .A(arr[605]), .B(n3470), .Y(n6163) );
  OAI21X1 U1246 ( .A(n5555), .B(n3466), .C(n6164), .Y(n8908) );
  NAND2X1 U1247 ( .A(arr[606]), .B(n3470), .Y(n6164) );
  OAI21X1 U1248 ( .A(n5557), .B(n3466), .C(n6165), .Y(n8909) );
  NAND2X1 U1249 ( .A(arr[607]), .B(n3470), .Y(n6165) );
  OAI21X1 U1250 ( .A(n5559), .B(n3465), .C(n6166), .Y(n8910) );
  NAND2X1 U1251 ( .A(arr[608]), .B(n3470), .Y(n6166) );
  OAI21X1 U1252 ( .A(n5561), .B(n3465), .C(n6167), .Y(n8911) );
  NAND2X1 U1253 ( .A(arr[609]), .B(n3470), .Y(n6167) );
  OAI21X1 U1254 ( .A(n5563), .B(n3465), .C(n6168), .Y(n8912) );
  NAND2X1 U1255 ( .A(arr[610]), .B(n3470), .Y(n6168) );
  OAI21X1 U1256 ( .A(n5565), .B(n3465), .C(n6169), .Y(n8913) );
  NAND2X1 U1257 ( .A(arr[611]), .B(n3470), .Y(n6169) );
  OAI21X1 U1258 ( .A(n5567), .B(n3465), .C(n6170), .Y(n8914) );
  NAND2X1 U1259 ( .A(arr[612]), .B(n3470), .Y(n6170) );
  OAI21X1 U1260 ( .A(n5569), .B(n3465), .C(n6171), .Y(n8915) );
  NAND2X1 U1261 ( .A(arr[613]), .B(n3468), .Y(n6171) );
  OAI21X1 U1262 ( .A(n5571), .B(n3465), .C(n6172), .Y(n8916) );
  NAND2X1 U1263 ( .A(arr[614]), .B(n3468), .Y(n6172) );
  NAND2X1 U1264 ( .A(n6088), .B(n5660), .Y(n6131) );
  OAI21X1 U1265 ( .A(n5491), .B(n3459), .C(n6174), .Y(n8917) );
  NAND2X1 U1266 ( .A(arr[615]), .B(n3462), .Y(n6174) );
  OAI21X1 U1267 ( .A(n5493), .B(n3459), .C(n6175), .Y(n8918) );
  NAND2X1 U1268 ( .A(arr[616]), .B(n3462), .Y(n6175) );
  OAI21X1 U1269 ( .A(n5495), .B(n3459), .C(n6176), .Y(n8919) );
  NAND2X1 U1270 ( .A(arr[617]), .B(n3462), .Y(n6176) );
  OAI21X1 U1271 ( .A(n5497), .B(n3459), .C(n6177), .Y(n8920) );
  NAND2X1 U1272 ( .A(arr[618]), .B(n3462), .Y(n6177) );
  OAI21X1 U1273 ( .A(n5499), .B(n3459), .C(n6178), .Y(n8921) );
  NAND2X1 U1274 ( .A(arr[619]), .B(n3462), .Y(n6178) );
  OAI21X1 U1275 ( .A(n5501), .B(n3460), .C(n6179), .Y(n8922) );
  NAND2X1 U1276 ( .A(arr[620]), .B(n3462), .Y(n6179) );
  OAI21X1 U1277 ( .A(n5503), .B(n3460), .C(n6180), .Y(n8923) );
  NAND2X1 U1278 ( .A(arr[621]), .B(n3462), .Y(n6180) );
  OAI21X1 U1279 ( .A(n5505), .B(n3460), .C(n6181), .Y(n8924) );
  NAND2X1 U1280 ( .A(arr[622]), .B(n3462), .Y(n6181) );
  OAI21X1 U1281 ( .A(n5507), .B(n3459), .C(n6182), .Y(n8925) );
  NAND2X1 U1282 ( .A(arr[623]), .B(n3462), .Y(n6182) );
  OAI21X1 U1283 ( .A(n5509), .B(n3460), .C(n6183), .Y(n8926) );
  NAND2X1 U1284 ( .A(arr[624]), .B(n3462), .Y(n6183) );
  OAI21X1 U1285 ( .A(n5511), .B(n3461), .C(n6184), .Y(n8927) );
  NAND2X1 U1286 ( .A(arr[625]), .B(n3462), .Y(n6184) );
  OAI21X1 U1287 ( .A(n5513), .B(n3461), .C(n6185), .Y(n8928) );
  NAND2X1 U1288 ( .A(arr[626]), .B(n3462), .Y(n6185) );
  OAI21X1 U1289 ( .A(n5515), .B(n3461), .C(n6186), .Y(n8929) );
  NAND2X1 U1290 ( .A(arr[627]), .B(n3462), .Y(n6186) );
  OAI21X1 U1291 ( .A(n5517), .B(n3460), .C(n6187), .Y(n8930) );
  NAND2X1 U1292 ( .A(arr[628]), .B(n3463), .Y(n6187) );
  OAI21X1 U1293 ( .A(n5519), .B(n3462), .C(n6188), .Y(n8931) );
  NAND2X1 U1294 ( .A(arr[629]), .B(n3463), .Y(n6188) );
  OAI21X1 U1295 ( .A(n5521), .B(n3462), .C(n6189), .Y(n8932) );
  NAND2X1 U1296 ( .A(arr[630]), .B(n3463), .Y(n6189) );
  OAI21X1 U1297 ( .A(n5523), .B(n3461), .C(n6190), .Y(n8933) );
  NAND2X1 U1298 ( .A(arr[631]), .B(n3463), .Y(n6190) );
  OAI21X1 U1299 ( .A(n5525), .B(n3461), .C(n6191), .Y(n8934) );
  NAND2X1 U1300 ( .A(arr[632]), .B(n3463), .Y(n6191) );
  OAI21X1 U1301 ( .A(n5527), .B(n3461), .C(n6192), .Y(n8935) );
  NAND2X1 U1302 ( .A(arr[633]), .B(n3463), .Y(n6192) );
  OAI21X1 U1303 ( .A(n5529), .B(n3461), .C(n6193), .Y(n8936) );
  NAND2X1 U1304 ( .A(arr[634]), .B(n3463), .Y(n6193) );
  OAI21X1 U1305 ( .A(n5531), .B(n3461), .C(n6194), .Y(n8937) );
  NAND2X1 U1306 ( .A(arr[635]), .B(n3463), .Y(n6194) );
  OAI21X1 U1307 ( .A(n5533), .B(n3461), .C(n6195), .Y(n8938) );
  NAND2X1 U1308 ( .A(arr[636]), .B(n3463), .Y(n6195) );
  OAI21X1 U1309 ( .A(n5535), .B(n3461), .C(n6196), .Y(n8939) );
  NAND2X1 U1310 ( .A(arr[637]), .B(n3463), .Y(n6196) );
  OAI21X1 U1311 ( .A(n5537), .B(n3461), .C(n6197), .Y(n8940) );
  NAND2X1 U1312 ( .A(arr[638]), .B(n3463), .Y(n6197) );
  OAI21X1 U1313 ( .A(n5539), .B(n3461), .C(n6198), .Y(n8941) );
  NAND2X1 U1314 ( .A(arr[639]), .B(n3463), .Y(n6198) );
  OAI21X1 U1315 ( .A(n5541), .B(n3461), .C(n6199), .Y(n8942) );
  NAND2X1 U1316 ( .A(arr[640]), .B(n3463), .Y(n6199) );
  OAI21X1 U1317 ( .A(n5543), .B(n3460), .C(n6200), .Y(n8943) );
  NAND2X1 U1318 ( .A(arr[641]), .B(n3463), .Y(n6200) );
  OAI21X1 U1319 ( .A(n5545), .B(n3460), .C(n6201), .Y(n8944) );
  NAND2X1 U1320 ( .A(arr[642]), .B(n3463), .Y(n6201) );
  OAI21X1 U1321 ( .A(n5547), .B(n3460), .C(n6202), .Y(n8945) );
  NAND2X1 U1322 ( .A(arr[643]), .B(n3463), .Y(n6202) );
  OAI21X1 U1323 ( .A(n5549), .B(n3460), .C(n6203), .Y(n8946) );
  NAND2X1 U1324 ( .A(arr[644]), .B(n3463), .Y(n6203) );
  OAI21X1 U1325 ( .A(n5551), .B(n3460), .C(n6204), .Y(n8947) );
  NAND2X1 U1326 ( .A(arr[645]), .B(n3464), .Y(n6204) );
  OAI21X1 U1327 ( .A(n5553), .B(n3460), .C(n6205), .Y(n8948) );
  NAND2X1 U1328 ( .A(arr[646]), .B(n3464), .Y(n6205) );
  OAI21X1 U1329 ( .A(n5555), .B(n3460), .C(n6206), .Y(n8949) );
  NAND2X1 U1330 ( .A(arr[647]), .B(n3464), .Y(n6206) );
  OAI21X1 U1331 ( .A(n5557), .B(n3460), .C(n6207), .Y(n8950) );
  NAND2X1 U1332 ( .A(arr[648]), .B(n3464), .Y(n6207) );
  OAI21X1 U1333 ( .A(n5559), .B(n3459), .C(n6208), .Y(n8951) );
  NAND2X1 U1334 ( .A(arr[649]), .B(n3464), .Y(n6208) );
  OAI21X1 U1335 ( .A(n5561), .B(n3459), .C(n6209), .Y(n8952) );
  NAND2X1 U1336 ( .A(arr[650]), .B(n3464), .Y(n6209) );
  OAI21X1 U1337 ( .A(n5563), .B(n3459), .C(n6210), .Y(n8953) );
  NAND2X1 U1338 ( .A(arr[651]), .B(n3464), .Y(n6210) );
  OAI21X1 U1339 ( .A(n5565), .B(n3459), .C(n6211), .Y(n8954) );
  NAND2X1 U1340 ( .A(arr[652]), .B(n3464), .Y(n6211) );
  OAI21X1 U1341 ( .A(n5567), .B(n3459), .C(n6212), .Y(n8955) );
  NAND2X1 U1342 ( .A(arr[653]), .B(n3464), .Y(n6212) );
  OAI21X1 U1343 ( .A(n5569), .B(n3459), .C(n6213), .Y(n8956) );
  NAND2X1 U1344 ( .A(arr[654]), .B(n3462), .Y(n6213) );
  OAI21X1 U1345 ( .A(n5571), .B(n3459), .C(n6214), .Y(n8957) );
  NAND2X1 U1346 ( .A(arr[655]), .B(n3462), .Y(n6214) );
  NAND2X1 U1347 ( .A(n6088), .B(n5703), .Y(n6173) );
  AND2X1 U1349 ( .A(n6216), .B(n6217), .Y(n5704) );
  OAI21X1 U1350 ( .A(n5491), .B(n3453), .C(n6219), .Y(n8958) );
  NAND2X1 U1351 ( .A(arr[656]), .B(n3456), .Y(n6219) );
  OAI21X1 U1352 ( .A(n5493), .B(n3453), .C(n6220), .Y(n8959) );
  NAND2X1 U1353 ( .A(arr[657]), .B(n3456), .Y(n6220) );
  OAI21X1 U1354 ( .A(n5495), .B(n3453), .C(n6221), .Y(n8960) );
  NAND2X1 U1355 ( .A(arr[658]), .B(n3456), .Y(n6221) );
  OAI21X1 U1356 ( .A(n5497), .B(n3453), .C(n6222), .Y(n8961) );
  NAND2X1 U1357 ( .A(arr[659]), .B(n3456), .Y(n6222) );
  OAI21X1 U1358 ( .A(n5499), .B(n3453), .C(n6223), .Y(n8962) );
  NAND2X1 U1359 ( .A(arr[660]), .B(n3456), .Y(n6223) );
  OAI21X1 U1360 ( .A(n5501), .B(n3454), .C(n6224), .Y(n8963) );
  NAND2X1 U1361 ( .A(arr[661]), .B(n3456), .Y(n6224) );
  OAI21X1 U1362 ( .A(n5503), .B(n3454), .C(n6225), .Y(n8964) );
  NAND2X1 U1363 ( .A(arr[662]), .B(n3456), .Y(n6225) );
  OAI21X1 U1364 ( .A(n5505), .B(n3454), .C(n6226), .Y(n8965) );
  NAND2X1 U1365 ( .A(arr[663]), .B(n3456), .Y(n6226) );
  OAI21X1 U1366 ( .A(n5507), .B(n3453), .C(n6227), .Y(n8966) );
  NAND2X1 U1367 ( .A(arr[664]), .B(n3456), .Y(n6227) );
  OAI21X1 U1368 ( .A(n5509), .B(n3454), .C(n6228), .Y(n8967) );
  NAND2X1 U1369 ( .A(arr[665]), .B(n3456), .Y(n6228) );
  OAI21X1 U1370 ( .A(n5511), .B(n3455), .C(n6229), .Y(n8968) );
  NAND2X1 U1371 ( .A(arr[666]), .B(n3456), .Y(n6229) );
  OAI21X1 U1372 ( .A(n5513), .B(n3455), .C(n6230), .Y(n8969) );
  NAND2X1 U1373 ( .A(arr[667]), .B(n3456), .Y(n6230) );
  OAI21X1 U1374 ( .A(n5515), .B(n3455), .C(n6231), .Y(n8970) );
  NAND2X1 U1375 ( .A(arr[668]), .B(n3456), .Y(n6231) );
  OAI21X1 U1376 ( .A(n5517), .B(n3454), .C(n6232), .Y(n8971) );
  NAND2X1 U1377 ( .A(arr[669]), .B(n3457), .Y(n6232) );
  OAI21X1 U1378 ( .A(n5519), .B(n3456), .C(n6233), .Y(n8972) );
  NAND2X1 U1379 ( .A(arr[670]), .B(n3457), .Y(n6233) );
  OAI21X1 U1380 ( .A(n5521), .B(n3456), .C(n6234), .Y(n8973) );
  NAND2X1 U1381 ( .A(arr[671]), .B(n3457), .Y(n6234) );
  OAI21X1 U1382 ( .A(n5523), .B(n3455), .C(n6235), .Y(n8974) );
  NAND2X1 U1383 ( .A(arr[672]), .B(n3457), .Y(n6235) );
  OAI21X1 U1384 ( .A(n5525), .B(n3455), .C(n6236), .Y(n8975) );
  NAND2X1 U1385 ( .A(arr[673]), .B(n3457), .Y(n6236) );
  OAI21X1 U1386 ( .A(n5527), .B(n3455), .C(n6237), .Y(n8976) );
  NAND2X1 U1387 ( .A(arr[674]), .B(n3457), .Y(n6237) );
  OAI21X1 U1388 ( .A(n5529), .B(n3455), .C(n6238), .Y(n8977) );
  NAND2X1 U1389 ( .A(arr[675]), .B(n3457), .Y(n6238) );
  OAI21X1 U1390 ( .A(n5531), .B(n3455), .C(n6239), .Y(n8978) );
  NAND2X1 U1391 ( .A(arr[676]), .B(n3457), .Y(n6239) );
  OAI21X1 U1392 ( .A(n5533), .B(n3455), .C(n6240), .Y(n8979) );
  NAND2X1 U1393 ( .A(arr[677]), .B(n3457), .Y(n6240) );
  OAI21X1 U1394 ( .A(n5535), .B(n3455), .C(n6241), .Y(n8980) );
  NAND2X1 U1395 ( .A(arr[678]), .B(n3457), .Y(n6241) );
  OAI21X1 U1396 ( .A(n5537), .B(n3455), .C(n6242), .Y(n8981) );
  NAND2X1 U1397 ( .A(arr[679]), .B(n3457), .Y(n6242) );
  OAI21X1 U1398 ( .A(n5539), .B(n3455), .C(n6243), .Y(n8982) );
  NAND2X1 U1399 ( .A(arr[680]), .B(n3457), .Y(n6243) );
  OAI21X1 U1400 ( .A(n5541), .B(n3455), .C(n6244), .Y(n8983) );
  NAND2X1 U1401 ( .A(arr[681]), .B(n3457), .Y(n6244) );
  OAI21X1 U1402 ( .A(n5543), .B(n3454), .C(n6245), .Y(n8984) );
  NAND2X1 U1403 ( .A(arr[682]), .B(n3457), .Y(n6245) );
  OAI21X1 U1404 ( .A(n5545), .B(n3454), .C(n6246), .Y(n8985) );
  NAND2X1 U1405 ( .A(arr[683]), .B(n3457), .Y(n6246) );
  OAI21X1 U1406 ( .A(n5547), .B(n3454), .C(n6247), .Y(n8986) );
  NAND2X1 U1407 ( .A(arr[684]), .B(n3457), .Y(n6247) );
  OAI21X1 U1408 ( .A(n5549), .B(n3454), .C(n6248), .Y(n8987) );
  NAND2X1 U1409 ( .A(arr[685]), .B(n3457), .Y(n6248) );
  OAI21X1 U1410 ( .A(n5551), .B(n3454), .C(n6249), .Y(n8988) );
  NAND2X1 U1411 ( .A(arr[686]), .B(n3458), .Y(n6249) );
  OAI21X1 U1412 ( .A(n5553), .B(n3454), .C(n6250), .Y(n8989) );
  NAND2X1 U1413 ( .A(arr[687]), .B(n3458), .Y(n6250) );
  OAI21X1 U1414 ( .A(n5555), .B(n3454), .C(n6251), .Y(n8990) );
  NAND2X1 U1415 ( .A(arr[688]), .B(n3458), .Y(n6251) );
  OAI21X1 U1416 ( .A(n5557), .B(n3454), .C(n6252), .Y(n8991) );
  NAND2X1 U1417 ( .A(arr[689]), .B(n3458), .Y(n6252) );
  OAI21X1 U1418 ( .A(n5559), .B(n3453), .C(n6253), .Y(n8992) );
  NAND2X1 U1419 ( .A(arr[690]), .B(n3458), .Y(n6253) );
  OAI21X1 U1420 ( .A(n5561), .B(n3453), .C(n6254), .Y(n8993) );
  NAND2X1 U1421 ( .A(arr[691]), .B(n3458), .Y(n6254) );
  OAI21X1 U1422 ( .A(n5563), .B(n3453), .C(n6255), .Y(n8994) );
  NAND2X1 U1423 ( .A(arr[692]), .B(n3458), .Y(n6255) );
  OAI21X1 U1424 ( .A(n5565), .B(n3453), .C(n6256), .Y(n8995) );
  NAND2X1 U1425 ( .A(arr[693]), .B(n3458), .Y(n6256) );
  OAI21X1 U1426 ( .A(n5567), .B(n3453), .C(n6257), .Y(n8996) );
  NAND2X1 U1427 ( .A(arr[694]), .B(n3458), .Y(n6257) );
  OAI21X1 U1428 ( .A(n5569), .B(n3453), .C(n6258), .Y(n8997) );
  NAND2X1 U1429 ( .A(arr[695]), .B(n3456), .Y(n6258) );
  OAI21X1 U1430 ( .A(n5571), .B(n3453), .C(n6259), .Y(n8998) );
  NAND2X1 U1431 ( .A(arr[696]), .B(n3456), .Y(n6259) );
  NAND2X1 U1432 ( .A(n6260), .B(n5573), .Y(n6218) );
  OAI21X1 U1433 ( .A(n5491), .B(n3447), .C(n6262), .Y(n8999) );
  NAND2X1 U1434 ( .A(arr[697]), .B(n3450), .Y(n6262) );
  OAI21X1 U1435 ( .A(n5493), .B(n3447), .C(n6263), .Y(n9000) );
  NAND2X1 U1436 ( .A(arr[698]), .B(n3450), .Y(n6263) );
  OAI21X1 U1437 ( .A(n5495), .B(n3447), .C(n6264), .Y(n9001) );
  NAND2X1 U1438 ( .A(arr[699]), .B(n3450), .Y(n6264) );
  OAI21X1 U1439 ( .A(n5497), .B(n3447), .C(n6265), .Y(n9002) );
  NAND2X1 U1440 ( .A(arr[700]), .B(n3450), .Y(n6265) );
  OAI21X1 U1441 ( .A(n5499), .B(n3447), .C(n6266), .Y(n9003) );
  NAND2X1 U1442 ( .A(arr[701]), .B(n3450), .Y(n6266) );
  OAI21X1 U1443 ( .A(n5501), .B(n3448), .C(n6267), .Y(n9004) );
  NAND2X1 U1444 ( .A(arr[702]), .B(n3450), .Y(n6267) );
  OAI21X1 U1445 ( .A(n5503), .B(n3448), .C(n6268), .Y(n9005) );
  NAND2X1 U1446 ( .A(arr[703]), .B(n3450), .Y(n6268) );
  OAI21X1 U1447 ( .A(n5505), .B(n3448), .C(n6269), .Y(n9006) );
  NAND2X1 U1448 ( .A(arr[704]), .B(n3450), .Y(n6269) );
  OAI21X1 U1449 ( .A(n5507), .B(n3447), .C(n6270), .Y(n9007) );
  NAND2X1 U1450 ( .A(arr[705]), .B(n3450), .Y(n6270) );
  OAI21X1 U1451 ( .A(n5509), .B(n3448), .C(n6271), .Y(n9008) );
  NAND2X1 U1452 ( .A(arr[706]), .B(n3450), .Y(n6271) );
  OAI21X1 U1453 ( .A(n5511), .B(n3449), .C(n6272), .Y(n9009) );
  NAND2X1 U1454 ( .A(arr[707]), .B(n3450), .Y(n6272) );
  OAI21X1 U1455 ( .A(n5513), .B(n3449), .C(n6273), .Y(n9010) );
  NAND2X1 U1456 ( .A(arr[708]), .B(n3450), .Y(n6273) );
  OAI21X1 U1457 ( .A(n5515), .B(n3449), .C(n6274), .Y(n9011) );
  NAND2X1 U1458 ( .A(arr[709]), .B(n3450), .Y(n6274) );
  OAI21X1 U1459 ( .A(n5517), .B(n3448), .C(n6275), .Y(n9012) );
  NAND2X1 U1460 ( .A(arr[710]), .B(n3451), .Y(n6275) );
  OAI21X1 U1461 ( .A(n5519), .B(n3450), .C(n6276), .Y(n9013) );
  NAND2X1 U1462 ( .A(arr[711]), .B(n3451), .Y(n6276) );
  OAI21X1 U1463 ( .A(n5521), .B(n3450), .C(n6277), .Y(n9014) );
  NAND2X1 U1464 ( .A(arr[712]), .B(n3451), .Y(n6277) );
  OAI21X1 U1465 ( .A(n5523), .B(n3449), .C(n6278), .Y(n9015) );
  NAND2X1 U1466 ( .A(arr[713]), .B(n3451), .Y(n6278) );
  OAI21X1 U1467 ( .A(n5525), .B(n3449), .C(n6279), .Y(n9016) );
  NAND2X1 U1468 ( .A(arr[714]), .B(n3451), .Y(n6279) );
  OAI21X1 U1469 ( .A(n5527), .B(n3449), .C(n6280), .Y(n9017) );
  NAND2X1 U1470 ( .A(arr[715]), .B(n3451), .Y(n6280) );
  OAI21X1 U1471 ( .A(n5529), .B(n3449), .C(n6281), .Y(n9018) );
  NAND2X1 U1472 ( .A(arr[716]), .B(n3451), .Y(n6281) );
  OAI21X1 U1473 ( .A(n5531), .B(n3449), .C(n6282), .Y(n9019) );
  NAND2X1 U1474 ( .A(arr[717]), .B(n3451), .Y(n6282) );
  OAI21X1 U1475 ( .A(n5533), .B(n3449), .C(n6283), .Y(n9020) );
  NAND2X1 U1476 ( .A(arr[718]), .B(n3451), .Y(n6283) );
  OAI21X1 U1477 ( .A(n5535), .B(n3449), .C(n6284), .Y(n9021) );
  NAND2X1 U1478 ( .A(arr[719]), .B(n3451), .Y(n6284) );
  OAI21X1 U1479 ( .A(n5537), .B(n3449), .C(n6285), .Y(n9022) );
  NAND2X1 U1480 ( .A(arr[720]), .B(n3451), .Y(n6285) );
  OAI21X1 U1481 ( .A(n5539), .B(n3449), .C(n6286), .Y(n9023) );
  NAND2X1 U1482 ( .A(arr[721]), .B(n3451), .Y(n6286) );
  OAI21X1 U1483 ( .A(n5541), .B(n3449), .C(n6287), .Y(n9024) );
  NAND2X1 U1484 ( .A(arr[722]), .B(n3451), .Y(n6287) );
  OAI21X1 U1485 ( .A(n5543), .B(n3448), .C(n6288), .Y(n9025) );
  NAND2X1 U1486 ( .A(arr[723]), .B(n3451), .Y(n6288) );
  OAI21X1 U1487 ( .A(n5545), .B(n3448), .C(n6289), .Y(n9026) );
  NAND2X1 U1488 ( .A(arr[724]), .B(n3451), .Y(n6289) );
  OAI21X1 U1489 ( .A(n5547), .B(n3448), .C(n6290), .Y(n9027) );
  NAND2X1 U1490 ( .A(arr[725]), .B(n3451), .Y(n6290) );
  OAI21X1 U1491 ( .A(n5549), .B(n3448), .C(n6291), .Y(n9028) );
  NAND2X1 U1492 ( .A(arr[726]), .B(n3451), .Y(n6291) );
  OAI21X1 U1493 ( .A(n5551), .B(n3448), .C(n6292), .Y(n9029) );
  NAND2X1 U1494 ( .A(arr[727]), .B(n3452), .Y(n6292) );
  OAI21X1 U1495 ( .A(n5553), .B(n3448), .C(n6293), .Y(n9030) );
  NAND2X1 U1496 ( .A(arr[728]), .B(n3452), .Y(n6293) );
  OAI21X1 U1497 ( .A(n5555), .B(n3448), .C(n6294), .Y(n9031) );
  NAND2X1 U1498 ( .A(arr[729]), .B(n3452), .Y(n6294) );
  OAI21X1 U1499 ( .A(n5557), .B(n3448), .C(n6295), .Y(n9032) );
  NAND2X1 U1500 ( .A(arr[730]), .B(n3452), .Y(n6295) );
  OAI21X1 U1501 ( .A(n5559), .B(n3447), .C(n6296), .Y(n9033) );
  NAND2X1 U1502 ( .A(arr[731]), .B(n3452), .Y(n6296) );
  OAI21X1 U1503 ( .A(n5561), .B(n3447), .C(n6297), .Y(n9034) );
  NAND2X1 U1504 ( .A(arr[732]), .B(n3452), .Y(n6297) );
  OAI21X1 U1505 ( .A(n5563), .B(n3447), .C(n6298), .Y(n9035) );
  NAND2X1 U1506 ( .A(arr[733]), .B(n3452), .Y(n6298) );
  OAI21X1 U1507 ( .A(n5565), .B(n3447), .C(n6299), .Y(n9036) );
  NAND2X1 U1508 ( .A(arr[734]), .B(n3452), .Y(n6299) );
  OAI21X1 U1509 ( .A(n5567), .B(n3447), .C(n6300), .Y(n9037) );
  NAND2X1 U1510 ( .A(arr[735]), .B(n3452), .Y(n6300) );
  OAI21X1 U1511 ( .A(n5569), .B(n3447), .C(n6301), .Y(n9038) );
  NAND2X1 U1512 ( .A(arr[736]), .B(n3450), .Y(n6301) );
  OAI21X1 U1513 ( .A(n5571), .B(n3447), .C(n6302), .Y(n9039) );
  NAND2X1 U1514 ( .A(arr[737]), .B(n3450), .Y(n6302) );
  NAND2X1 U1515 ( .A(n6260), .B(n5617), .Y(n6261) );
  OAI21X1 U1516 ( .A(n5491), .B(n3441), .C(n6304), .Y(n9040) );
  NAND2X1 U1517 ( .A(arr[738]), .B(n3444), .Y(n6304) );
  OAI21X1 U1518 ( .A(n5493), .B(n3441), .C(n6305), .Y(n9041) );
  NAND2X1 U1519 ( .A(arr[739]), .B(n3444), .Y(n6305) );
  OAI21X1 U1520 ( .A(n5495), .B(n3441), .C(n6306), .Y(n9042) );
  NAND2X1 U1521 ( .A(arr[740]), .B(n3444), .Y(n6306) );
  OAI21X1 U1522 ( .A(n5497), .B(n3441), .C(n6307), .Y(n9043) );
  NAND2X1 U1523 ( .A(arr[741]), .B(n3444), .Y(n6307) );
  OAI21X1 U1524 ( .A(n5499), .B(n3441), .C(n6308), .Y(n9044) );
  NAND2X1 U1525 ( .A(arr[742]), .B(n3444), .Y(n6308) );
  OAI21X1 U1526 ( .A(n5501), .B(n3442), .C(n6309), .Y(n9045) );
  NAND2X1 U1527 ( .A(arr[743]), .B(n3444), .Y(n6309) );
  OAI21X1 U1528 ( .A(n5503), .B(n3442), .C(n6310), .Y(n9046) );
  NAND2X1 U1529 ( .A(arr[744]), .B(n3444), .Y(n6310) );
  OAI21X1 U1530 ( .A(n5505), .B(n3442), .C(n6311), .Y(n9047) );
  NAND2X1 U1531 ( .A(arr[745]), .B(n3444), .Y(n6311) );
  OAI21X1 U1532 ( .A(n5507), .B(n3441), .C(n6312), .Y(n9048) );
  NAND2X1 U1533 ( .A(arr[746]), .B(n3444), .Y(n6312) );
  OAI21X1 U1534 ( .A(n5509), .B(n3442), .C(n6313), .Y(n9049) );
  NAND2X1 U1535 ( .A(arr[747]), .B(n3444), .Y(n6313) );
  OAI21X1 U1536 ( .A(n5511), .B(n3443), .C(n6314), .Y(n9050) );
  NAND2X1 U1537 ( .A(arr[748]), .B(n3444), .Y(n6314) );
  OAI21X1 U1538 ( .A(n5513), .B(n3443), .C(n6315), .Y(n9051) );
  NAND2X1 U1539 ( .A(arr[749]), .B(n3444), .Y(n6315) );
  OAI21X1 U1540 ( .A(n5515), .B(n3443), .C(n6316), .Y(n9052) );
  NAND2X1 U1541 ( .A(arr[750]), .B(n3444), .Y(n6316) );
  OAI21X1 U1542 ( .A(n5517), .B(n3442), .C(n6317), .Y(n9053) );
  NAND2X1 U1543 ( .A(arr[751]), .B(n3445), .Y(n6317) );
  OAI21X1 U1544 ( .A(n5519), .B(n3444), .C(n6318), .Y(n9054) );
  NAND2X1 U1545 ( .A(arr[752]), .B(n3445), .Y(n6318) );
  OAI21X1 U1546 ( .A(n5521), .B(n3444), .C(n6319), .Y(n9055) );
  NAND2X1 U1547 ( .A(arr[753]), .B(n3445), .Y(n6319) );
  OAI21X1 U1548 ( .A(n5523), .B(n3443), .C(n6320), .Y(n9056) );
  NAND2X1 U1549 ( .A(arr[754]), .B(n3445), .Y(n6320) );
  OAI21X1 U1550 ( .A(n5525), .B(n3443), .C(n6321), .Y(n9057) );
  NAND2X1 U1551 ( .A(arr[755]), .B(n3445), .Y(n6321) );
  OAI21X1 U1552 ( .A(n5527), .B(n3443), .C(n6322), .Y(n9058) );
  NAND2X1 U1553 ( .A(arr[756]), .B(n3445), .Y(n6322) );
  OAI21X1 U1554 ( .A(n5529), .B(n3443), .C(n6323), .Y(n9059) );
  NAND2X1 U1555 ( .A(arr[757]), .B(n3445), .Y(n6323) );
  OAI21X1 U1556 ( .A(n5531), .B(n3443), .C(n6324), .Y(n9060) );
  NAND2X1 U1557 ( .A(arr[758]), .B(n3445), .Y(n6324) );
  OAI21X1 U1558 ( .A(n5533), .B(n3443), .C(n6325), .Y(n9061) );
  NAND2X1 U1559 ( .A(arr[759]), .B(n3445), .Y(n6325) );
  OAI21X1 U1560 ( .A(n5535), .B(n3443), .C(n6326), .Y(n9062) );
  NAND2X1 U1561 ( .A(arr[760]), .B(n3445), .Y(n6326) );
  OAI21X1 U1562 ( .A(n5537), .B(n3443), .C(n6327), .Y(n9063) );
  NAND2X1 U1563 ( .A(arr[761]), .B(n3445), .Y(n6327) );
  OAI21X1 U1564 ( .A(n5539), .B(n3443), .C(n6328), .Y(n9064) );
  NAND2X1 U1565 ( .A(arr[762]), .B(n3445), .Y(n6328) );
  OAI21X1 U1566 ( .A(n5541), .B(n3443), .C(n6329), .Y(n9065) );
  NAND2X1 U1567 ( .A(arr[763]), .B(n3445), .Y(n6329) );
  OAI21X1 U1568 ( .A(n5543), .B(n3442), .C(n6330), .Y(n9066) );
  NAND2X1 U1569 ( .A(arr[764]), .B(n3445), .Y(n6330) );
  OAI21X1 U1570 ( .A(n5545), .B(n3442), .C(n6331), .Y(n9067) );
  NAND2X1 U1571 ( .A(arr[765]), .B(n3445), .Y(n6331) );
  OAI21X1 U1572 ( .A(n5547), .B(n3442), .C(n6332), .Y(n9068) );
  NAND2X1 U1573 ( .A(arr[766]), .B(n3445), .Y(n6332) );
  OAI21X1 U1574 ( .A(n5549), .B(n3442), .C(n6333), .Y(n9069) );
  NAND2X1 U1575 ( .A(arr[767]), .B(n3445), .Y(n6333) );
  OAI21X1 U1576 ( .A(n5551), .B(n3442), .C(n6334), .Y(n9070) );
  NAND2X1 U1577 ( .A(arr[768]), .B(n3446), .Y(n6334) );
  OAI21X1 U1578 ( .A(n5553), .B(n3442), .C(n6335), .Y(n9071) );
  NAND2X1 U1579 ( .A(arr[769]), .B(n3446), .Y(n6335) );
  OAI21X1 U1580 ( .A(n5555), .B(n3442), .C(n6336), .Y(n9072) );
  NAND2X1 U1581 ( .A(arr[770]), .B(n3446), .Y(n6336) );
  OAI21X1 U1582 ( .A(n5557), .B(n3442), .C(n6337), .Y(n9073) );
  NAND2X1 U1583 ( .A(arr[771]), .B(n3446), .Y(n6337) );
  OAI21X1 U1584 ( .A(n5559), .B(n3441), .C(n6338), .Y(n9074) );
  NAND2X1 U1585 ( .A(arr[772]), .B(n3446), .Y(n6338) );
  OAI21X1 U1586 ( .A(n5561), .B(n3441), .C(n6339), .Y(n9075) );
  NAND2X1 U1587 ( .A(arr[773]), .B(n3446), .Y(n6339) );
  OAI21X1 U1588 ( .A(n5563), .B(n3441), .C(n6340), .Y(n9076) );
  NAND2X1 U1589 ( .A(arr[774]), .B(n3446), .Y(n6340) );
  OAI21X1 U1590 ( .A(n5565), .B(n3441), .C(n6341), .Y(n9077) );
  NAND2X1 U1591 ( .A(arr[775]), .B(n3446), .Y(n6341) );
  OAI21X1 U1592 ( .A(n5567), .B(n3441), .C(n6342), .Y(n9078) );
  NAND2X1 U1593 ( .A(arr[776]), .B(n3446), .Y(n6342) );
  OAI21X1 U1594 ( .A(n5569), .B(n3441), .C(n6343), .Y(n9079) );
  NAND2X1 U1595 ( .A(arr[777]), .B(n3444), .Y(n6343) );
  OAI21X1 U1596 ( .A(n5571), .B(n3441), .C(n6344), .Y(n9080) );
  NAND2X1 U1597 ( .A(arr[778]), .B(n3444), .Y(n6344) );
  NAND2X1 U1598 ( .A(n6260), .B(n5660), .Y(n6303) );
  OAI21X1 U1599 ( .A(n5491), .B(n3435), .C(n6346), .Y(n9081) );
  NAND2X1 U1600 ( .A(arr[779]), .B(n3438), .Y(n6346) );
  OAI21X1 U1601 ( .A(n5493), .B(n3435), .C(n6347), .Y(n9082) );
  NAND2X1 U1602 ( .A(arr[780]), .B(n3438), .Y(n6347) );
  OAI21X1 U1603 ( .A(n5495), .B(n3435), .C(n6348), .Y(n9083) );
  NAND2X1 U1604 ( .A(arr[781]), .B(n3438), .Y(n6348) );
  OAI21X1 U1605 ( .A(n5497), .B(n3435), .C(n6349), .Y(n9084) );
  NAND2X1 U1606 ( .A(arr[782]), .B(n3438), .Y(n6349) );
  OAI21X1 U1607 ( .A(n5499), .B(n3435), .C(n6350), .Y(n9085) );
  NAND2X1 U1608 ( .A(arr[783]), .B(n3438), .Y(n6350) );
  OAI21X1 U1609 ( .A(n5501), .B(n3436), .C(n6351), .Y(n9086) );
  NAND2X1 U1610 ( .A(arr[784]), .B(n3438), .Y(n6351) );
  OAI21X1 U1611 ( .A(n5503), .B(n3436), .C(n6352), .Y(n9087) );
  NAND2X1 U1612 ( .A(arr[785]), .B(n3438), .Y(n6352) );
  OAI21X1 U1613 ( .A(n5505), .B(n3436), .C(n6353), .Y(n9088) );
  NAND2X1 U1614 ( .A(arr[786]), .B(n3438), .Y(n6353) );
  OAI21X1 U1615 ( .A(n5507), .B(n3435), .C(n6354), .Y(n9089) );
  NAND2X1 U1616 ( .A(arr[787]), .B(n3438), .Y(n6354) );
  OAI21X1 U1617 ( .A(n5509), .B(n3436), .C(n6355), .Y(n9090) );
  NAND2X1 U1618 ( .A(arr[788]), .B(n3438), .Y(n6355) );
  OAI21X1 U1619 ( .A(n5511), .B(n3437), .C(n6356), .Y(n9091) );
  NAND2X1 U1620 ( .A(arr[789]), .B(n3438), .Y(n6356) );
  OAI21X1 U1621 ( .A(n5513), .B(n3437), .C(n6357), .Y(n9092) );
  NAND2X1 U1622 ( .A(arr[790]), .B(n3438), .Y(n6357) );
  OAI21X1 U1623 ( .A(n5515), .B(n3437), .C(n6358), .Y(n9093) );
  NAND2X1 U1624 ( .A(arr[791]), .B(n3438), .Y(n6358) );
  OAI21X1 U1625 ( .A(n5517), .B(n3436), .C(n6359), .Y(n9094) );
  NAND2X1 U1626 ( .A(arr[792]), .B(n3439), .Y(n6359) );
  OAI21X1 U1627 ( .A(n5519), .B(n3438), .C(n6360), .Y(n9095) );
  NAND2X1 U1628 ( .A(arr[793]), .B(n3439), .Y(n6360) );
  OAI21X1 U1629 ( .A(n5521), .B(n3438), .C(n6361), .Y(n9096) );
  NAND2X1 U1630 ( .A(arr[794]), .B(n3439), .Y(n6361) );
  OAI21X1 U1631 ( .A(n5523), .B(n3437), .C(n6362), .Y(n9097) );
  NAND2X1 U1632 ( .A(arr[795]), .B(n3439), .Y(n6362) );
  OAI21X1 U1633 ( .A(n5525), .B(n3437), .C(n6363), .Y(n9098) );
  NAND2X1 U1634 ( .A(arr[796]), .B(n3439), .Y(n6363) );
  OAI21X1 U1635 ( .A(n5527), .B(n3437), .C(n6364), .Y(n9099) );
  NAND2X1 U1636 ( .A(arr[797]), .B(n3439), .Y(n6364) );
  OAI21X1 U1637 ( .A(n5529), .B(n3437), .C(n6365), .Y(n9100) );
  NAND2X1 U1638 ( .A(arr[798]), .B(n3439), .Y(n6365) );
  OAI21X1 U1639 ( .A(n5531), .B(n3437), .C(n6366), .Y(n9101) );
  NAND2X1 U1640 ( .A(arr[799]), .B(n3439), .Y(n6366) );
  OAI21X1 U1641 ( .A(n5533), .B(n3437), .C(n6367), .Y(n9102) );
  NAND2X1 U1642 ( .A(arr[800]), .B(n3439), .Y(n6367) );
  OAI21X1 U1643 ( .A(n5535), .B(n3437), .C(n6368), .Y(n9103) );
  NAND2X1 U1644 ( .A(arr[801]), .B(n3439), .Y(n6368) );
  OAI21X1 U1645 ( .A(n5537), .B(n3437), .C(n6369), .Y(n9104) );
  NAND2X1 U1646 ( .A(arr[802]), .B(n3439), .Y(n6369) );
  OAI21X1 U1647 ( .A(n5539), .B(n3437), .C(n6370), .Y(n9105) );
  NAND2X1 U1648 ( .A(arr[803]), .B(n3439), .Y(n6370) );
  OAI21X1 U1649 ( .A(n5541), .B(n3437), .C(n6371), .Y(n9106) );
  NAND2X1 U1650 ( .A(arr[804]), .B(n3439), .Y(n6371) );
  OAI21X1 U1651 ( .A(n5543), .B(n3436), .C(n6372), .Y(n9107) );
  NAND2X1 U1652 ( .A(arr[805]), .B(n3439), .Y(n6372) );
  OAI21X1 U1653 ( .A(n5545), .B(n3436), .C(n6373), .Y(n9108) );
  NAND2X1 U1654 ( .A(arr[806]), .B(n3439), .Y(n6373) );
  OAI21X1 U1655 ( .A(n5547), .B(n3436), .C(n6374), .Y(n9109) );
  NAND2X1 U1656 ( .A(arr[807]), .B(n3439), .Y(n6374) );
  OAI21X1 U1657 ( .A(n5549), .B(n3436), .C(n6375), .Y(n9110) );
  NAND2X1 U1658 ( .A(arr[808]), .B(n3439), .Y(n6375) );
  OAI21X1 U1659 ( .A(n5551), .B(n3436), .C(n6376), .Y(n9111) );
  NAND2X1 U1660 ( .A(arr[809]), .B(n3440), .Y(n6376) );
  OAI21X1 U1661 ( .A(n5553), .B(n3436), .C(n6377), .Y(n9112) );
  NAND2X1 U1662 ( .A(arr[810]), .B(n3440), .Y(n6377) );
  OAI21X1 U1663 ( .A(n5555), .B(n3436), .C(n6378), .Y(n9113) );
  NAND2X1 U1664 ( .A(arr[811]), .B(n3440), .Y(n6378) );
  OAI21X1 U1665 ( .A(n5557), .B(n3436), .C(n6379), .Y(n9114) );
  NAND2X1 U1666 ( .A(arr[812]), .B(n3440), .Y(n6379) );
  OAI21X1 U1667 ( .A(n5559), .B(n3435), .C(n6380), .Y(n9115) );
  NAND2X1 U1668 ( .A(arr[813]), .B(n3440), .Y(n6380) );
  OAI21X1 U1669 ( .A(n5561), .B(n3435), .C(n6381), .Y(n9116) );
  NAND2X1 U1670 ( .A(arr[814]), .B(n3440), .Y(n6381) );
  OAI21X1 U1671 ( .A(n5563), .B(n3435), .C(n6382), .Y(n9117) );
  NAND2X1 U1672 ( .A(arr[815]), .B(n3440), .Y(n6382) );
  OAI21X1 U1673 ( .A(n5565), .B(n3435), .C(n6383), .Y(n9118) );
  NAND2X1 U1674 ( .A(arr[816]), .B(n3440), .Y(n6383) );
  OAI21X1 U1675 ( .A(n5567), .B(n3435), .C(n6384), .Y(n9119) );
  NAND2X1 U1676 ( .A(arr[817]), .B(n3440), .Y(n6384) );
  OAI21X1 U1677 ( .A(n5569), .B(n3435), .C(n6385), .Y(n9120) );
  NAND2X1 U1678 ( .A(arr[818]), .B(n3438), .Y(n6385) );
  OAI21X1 U1679 ( .A(n5571), .B(n3435), .C(n6386), .Y(n9121) );
  NAND2X1 U1680 ( .A(arr[819]), .B(n3438), .Y(n6386) );
  NAND2X1 U1681 ( .A(n6260), .B(n5703), .Y(n6345) );
  OAI21X1 U1683 ( .A(n5491), .B(n3429), .C(n6389), .Y(n9122) );
  NAND2X1 U1684 ( .A(arr[820]), .B(n3432), .Y(n6389) );
  OAI21X1 U1685 ( .A(n5493), .B(n3429), .C(n6390), .Y(n9123) );
  NAND2X1 U1686 ( .A(arr[821]), .B(n3432), .Y(n6390) );
  OAI21X1 U1687 ( .A(n5495), .B(n3429), .C(n6391), .Y(n9124) );
  NAND2X1 U1688 ( .A(arr[822]), .B(n3432), .Y(n6391) );
  OAI21X1 U1689 ( .A(n5497), .B(n3429), .C(n6392), .Y(n9125) );
  NAND2X1 U1690 ( .A(arr[823]), .B(n3432), .Y(n6392) );
  OAI21X1 U1691 ( .A(n5499), .B(n3429), .C(n6393), .Y(n9126) );
  NAND2X1 U1692 ( .A(arr[824]), .B(n3432), .Y(n6393) );
  OAI21X1 U1693 ( .A(n5501), .B(n3430), .C(n6394), .Y(n9127) );
  NAND2X1 U1694 ( .A(arr[825]), .B(n3432), .Y(n6394) );
  OAI21X1 U1695 ( .A(n5503), .B(n3430), .C(n6395), .Y(n9128) );
  NAND2X1 U1696 ( .A(arr[826]), .B(n3432), .Y(n6395) );
  OAI21X1 U1697 ( .A(n5505), .B(n3430), .C(n6396), .Y(n9129) );
  NAND2X1 U1698 ( .A(arr[827]), .B(n3432), .Y(n6396) );
  OAI21X1 U1699 ( .A(n5507), .B(n3429), .C(n6397), .Y(n9130) );
  NAND2X1 U1700 ( .A(arr[828]), .B(n3432), .Y(n6397) );
  OAI21X1 U1701 ( .A(n5509), .B(n3430), .C(n6398), .Y(n9131) );
  NAND2X1 U1702 ( .A(arr[829]), .B(n3432), .Y(n6398) );
  OAI21X1 U1703 ( .A(n5511), .B(n3431), .C(n6399), .Y(n9132) );
  NAND2X1 U1704 ( .A(arr[830]), .B(n3432), .Y(n6399) );
  OAI21X1 U1705 ( .A(n5513), .B(n3431), .C(n6400), .Y(n9133) );
  NAND2X1 U1706 ( .A(arr[831]), .B(n3432), .Y(n6400) );
  OAI21X1 U1707 ( .A(n5515), .B(n3431), .C(n6401), .Y(n9134) );
  NAND2X1 U1708 ( .A(arr[832]), .B(n3432), .Y(n6401) );
  OAI21X1 U1709 ( .A(n5517), .B(n3430), .C(n6402), .Y(n9135) );
  NAND2X1 U1710 ( .A(arr[833]), .B(n3433), .Y(n6402) );
  OAI21X1 U1711 ( .A(n5519), .B(n3432), .C(n6403), .Y(n9136) );
  NAND2X1 U1712 ( .A(arr[834]), .B(n3433), .Y(n6403) );
  OAI21X1 U1713 ( .A(n5521), .B(n3432), .C(n6404), .Y(n9137) );
  NAND2X1 U1714 ( .A(arr[835]), .B(n3433), .Y(n6404) );
  OAI21X1 U1715 ( .A(n5523), .B(n3431), .C(n6405), .Y(n9138) );
  NAND2X1 U1716 ( .A(arr[836]), .B(n3433), .Y(n6405) );
  OAI21X1 U1717 ( .A(n5525), .B(n3431), .C(n6406), .Y(n9139) );
  NAND2X1 U1718 ( .A(arr[837]), .B(n3433), .Y(n6406) );
  OAI21X1 U1719 ( .A(n5527), .B(n3431), .C(n6407), .Y(n9140) );
  NAND2X1 U1720 ( .A(arr[838]), .B(n3433), .Y(n6407) );
  OAI21X1 U1721 ( .A(n5529), .B(n3431), .C(n6408), .Y(n9141) );
  NAND2X1 U1722 ( .A(arr[839]), .B(n3433), .Y(n6408) );
  OAI21X1 U1723 ( .A(n5531), .B(n3431), .C(n6409), .Y(n9142) );
  NAND2X1 U1724 ( .A(arr[840]), .B(n3433), .Y(n6409) );
  OAI21X1 U1725 ( .A(n5533), .B(n3431), .C(n6410), .Y(n9143) );
  NAND2X1 U1726 ( .A(arr[841]), .B(n3433), .Y(n6410) );
  OAI21X1 U1727 ( .A(n5535), .B(n3431), .C(n6411), .Y(n9144) );
  NAND2X1 U1728 ( .A(arr[842]), .B(n3433), .Y(n6411) );
  OAI21X1 U1729 ( .A(n5537), .B(n3431), .C(n6412), .Y(n9145) );
  NAND2X1 U1730 ( .A(arr[843]), .B(n3433), .Y(n6412) );
  OAI21X1 U1731 ( .A(n5539), .B(n3431), .C(n6413), .Y(n9146) );
  NAND2X1 U1732 ( .A(arr[844]), .B(n3433), .Y(n6413) );
  OAI21X1 U1733 ( .A(n5541), .B(n3431), .C(n6414), .Y(n9147) );
  NAND2X1 U1734 ( .A(arr[845]), .B(n3433), .Y(n6414) );
  OAI21X1 U1735 ( .A(n5543), .B(n3430), .C(n6415), .Y(n9148) );
  NAND2X1 U1736 ( .A(arr[846]), .B(n3433), .Y(n6415) );
  OAI21X1 U1737 ( .A(n5545), .B(n3430), .C(n6416), .Y(n9149) );
  NAND2X1 U1738 ( .A(arr[847]), .B(n3433), .Y(n6416) );
  OAI21X1 U1739 ( .A(n5547), .B(n3430), .C(n6417), .Y(n9150) );
  NAND2X1 U1740 ( .A(arr[848]), .B(n3433), .Y(n6417) );
  OAI21X1 U1741 ( .A(n5549), .B(n3430), .C(n6418), .Y(n9151) );
  NAND2X1 U1742 ( .A(arr[849]), .B(n3433), .Y(n6418) );
  OAI21X1 U1743 ( .A(n5551), .B(n3430), .C(n6419), .Y(n9152) );
  NAND2X1 U1744 ( .A(arr[850]), .B(n3434), .Y(n6419) );
  OAI21X1 U1745 ( .A(n5553), .B(n3430), .C(n6420), .Y(n9153) );
  NAND2X1 U1746 ( .A(arr[851]), .B(n3434), .Y(n6420) );
  OAI21X1 U1747 ( .A(n5555), .B(n3430), .C(n6421), .Y(n9154) );
  NAND2X1 U1748 ( .A(arr[852]), .B(n3434), .Y(n6421) );
  OAI21X1 U1749 ( .A(n5557), .B(n3430), .C(n6422), .Y(n9155) );
  NAND2X1 U1750 ( .A(arr[853]), .B(n3434), .Y(n6422) );
  OAI21X1 U1751 ( .A(n5559), .B(n3429), .C(n6423), .Y(n9156) );
  NAND2X1 U1752 ( .A(arr[854]), .B(n3434), .Y(n6423) );
  OAI21X1 U1753 ( .A(n5561), .B(n3429), .C(n6424), .Y(n9157) );
  NAND2X1 U1754 ( .A(arr[855]), .B(n3434), .Y(n6424) );
  OAI21X1 U1755 ( .A(n5563), .B(n3429), .C(n6425), .Y(n9158) );
  NAND2X1 U1756 ( .A(arr[856]), .B(n3434), .Y(n6425) );
  OAI21X1 U1757 ( .A(n5565), .B(n3429), .C(n6426), .Y(n9159) );
  NAND2X1 U1758 ( .A(arr[857]), .B(n3434), .Y(n6426) );
  OAI21X1 U1759 ( .A(n5567), .B(n3429), .C(n6427), .Y(n9160) );
  NAND2X1 U1760 ( .A(arr[858]), .B(n3434), .Y(n6427) );
  OAI21X1 U1761 ( .A(n5569), .B(n3429), .C(n6428), .Y(n9161) );
  NAND2X1 U1762 ( .A(arr[859]), .B(n3432), .Y(n6428) );
  OAI21X1 U1763 ( .A(n5571), .B(n3429), .C(n6429), .Y(n9162) );
  NAND2X1 U1764 ( .A(arr[860]), .B(n3432), .Y(n6429) );
  NAND2X1 U1765 ( .A(n6430), .B(n5573), .Y(n6388) );
  OAI21X1 U1766 ( .A(n5491), .B(n3423), .C(n6432), .Y(n9163) );
  NAND2X1 U1767 ( .A(arr[861]), .B(n3426), .Y(n6432) );
  OAI21X1 U1768 ( .A(n5493), .B(n3423), .C(n6433), .Y(n9164) );
  NAND2X1 U1769 ( .A(arr[862]), .B(n3426), .Y(n6433) );
  OAI21X1 U1770 ( .A(n5495), .B(n3423), .C(n6434), .Y(n9165) );
  NAND2X1 U1771 ( .A(arr[863]), .B(n3426), .Y(n6434) );
  OAI21X1 U1772 ( .A(n5497), .B(n3423), .C(n6435), .Y(n9166) );
  NAND2X1 U1773 ( .A(arr[864]), .B(n3426), .Y(n6435) );
  OAI21X1 U1774 ( .A(n5499), .B(n3423), .C(n6436), .Y(n9167) );
  NAND2X1 U1775 ( .A(arr[865]), .B(n3426), .Y(n6436) );
  OAI21X1 U1776 ( .A(n5501), .B(n3424), .C(n6437), .Y(n9168) );
  NAND2X1 U1777 ( .A(arr[866]), .B(n3426), .Y(n6437) );
  OAI21X1 U1778 ( .A(n5503), .B(n3424), .C(n6438), .Y(n9169) );
  NAND2X1 U1779 ( .A(arr[867]), .B(n3426), .Y(n6438) );
  OAI21X1 U1780 ( .A(n5505), .B(n3424), .C(n6439), .Y(n9170) );
  NAND2X1 U1781 ( .A(arr[868]), .B(n3426), .Y(n6439) );
  OAI21X1 U1782 ( .A(n5507), .B(n3423), .C(n6440), .Y(n9171) );
  NAND2X1 U1783 ( .A(arr[869]), .B(n3426), .Y(n6440) );
  OAI21X1 U1784 ( .A(n5509), .B(n3424), .C(n6441), .Y(n9172) );
  NAND2X1 U1785 ( .A(arr[870]), .B(n3426), .Y(n6441) );
  OAI21X1 U1786 ( .A(n5511), .B(n3425), .C(n6442), .Y(n9173) );
  NAND2X1 U1787 ( .A(arr[871]), .B(n3426), .Y(n6442) );
  OAI21X1 U1788 ( .A(n5513), .B(n3425), .C(n6443), .Y(n9174) );
  NAND2X1 U1789 ( .A(arr[872]), .B(n3426), .Y(n6443) );
  OAI21X1 U1790 ( .A(n5515), .B(n3425), .C(n6444), .Y(n9175) );
  NAND2X1 U1791 ( .A(arr[873]), .B(n3426), .Y(n6444) );
  OAI21X1 U1792 ( .A(n5517), .B(n3424), .C(n6445), .Y(n9176) );
  NAND2X1 U1793 ( .A(arr[874]), .B(n3427), .Y(n6445) );
  OAI21X1 U1794 ( .A(n5519), .B(n3426), .C(n6446), .Y(n9177) );
  NAND2X1 U1795 ( .A(arr[875]), .B(n3427), .Y(n6446) );
  OAI21X1 U1796 ( .A(n5521), .B(n3426), .C(n6447), .Y(n9178) );
  NAND2X1 U1797 ( .A(arr[876]), .B(n3427), .Y(n6447) );
  OAI21X1 U1798 ( .A(n5523), .B(n3425), .C(n6448), .Y(n9179) );
  NAND2X1 U1799 ( .A(arr[877]), .B(n3427), .Y(n6448) );
  OAI21X1 U1800 ( .A(n5525), .B(n3425), .C(n6449), .Y(n9180) );
  NAND2X1 U1801 ( .A(arr[878]), .B(n3427), .Y(n6449) );
  OAI21X1 U1802 ( .A(n5527), .B(n3425), .C(n6450), .Y(n9181) );
  NAND2X1 U1803 ( .A(arr[879]), .B(n3427), .Y(n6450) );
  OAI21X1 U1804 ( .A(n5529), .B(n3425), .C(n6451), .Y(n9182) );
  NAND2X1 U1805 ( .A(arr[880]), .B(n3427), .Y(n6451) );
  OAI21X1 U1806 ( .A(n5531), .B(n3425), .C(n6452), .Y(n9183) );
  NAND2X1 U1807 ( .A(arr[881]), .B(n3427), .Y(n6452) );
  OAI21X1 U1808 ( .A(n5533), .B(n3425), .C(n6453), .Y(n9184) );
  NAND2X1 U1809 ( .A(arr[882]), .B(n3427), .Y(n6453) );
  OAI21X1 U1810 ( .A(n5535), .B(n3425), .C(n6454), .Y(n9185) );
  NAND2X1 U1811 ( .A(arr[883]), .B(n3427), .Y(n6454) );
  OAI21X1 U1812 ( .A(n5537), .B(n3425), .C(n6455), .Y(n9186) );
  NAND2X1 U1813 ( .A(arr[884]), .B(n3427), .Y(n6455) );
  OAI21X1 U1814 ( .A(n5539), .B(n3425), .C(n6456), .Y(n9187) );
  NAND2X1 U1815 ( .A(arr[885]), .B(n3427), .Y(n6456) );
  OAI21X1 U1816 ( .A(n5541), .B(n3425), .C(n6457), .Y(n9188) );
  NAND2X1 U1817 ( .A(arr[886]), .B(n3427), .Y(n6457) );
  OAI21X1 U1818 ( .A(n5543), .B(n3424), .C(n6458), .Y(n9189) );
  NAND2X1 U1819 ( .A(arr[887]), .B(n3427), .Y(n6458) );
  OAI21X1 U1820 ( .A(n5545), .B(n3424), .C(n6459), .Y(n9190) );
  NAND2X1 U1821 ( .A(arr[888]), .B(n3427), .Y(n6459) );
  OAI21X1 U1822 ( .A(n5547), .B(n3424), .C(n6460), .Y(n9191) );
  NAND2X1 U1823 ( .A(arr[889]), .B(n3427), .Y(n6460) );
  OAI21X1 U1824 ( .A(n5549), .B(n3424), .C(n6461), .Y(n9192) );
  NAND2X1 U1825 ( .A(arr[890]), .B(n3427), .Y(n6461) );
  OAI21X1 U1826 ( .A(n5551), .B(n3424), .C(n6462), .Y(n9193) );
  NAND2X1 U1827 ( .A(arr[891]), .B(n3428), .Y(n6462) );
  OAI21X1 U1828 ( .A(n5553), .B(n3424), .C(n6463), .Y(n9194) );
  NAND2X1 U1829 ( .A(arr[892]), .B(n3428), .Y(n6463) );
  OAI21X1 U1830 ( .A(n5555), .B(n3424), .C(n6464), .Y(n9195) );
  NAND2X1 U1831 ( .A(arr[893]), .B(n3428), .Y(n6464) );
  OAI21X1 U1832 ( .A(n5557), .B(n3424), .C(n6465), .Y(n9196) );
  NAND2X1 U1833 ( .A(arr[894]), .B(n3428), .Y(n6465) );
  OAI21X1 U1834 ( .A(n5559), .B(n3423), .C(n6466), .Y(n9197) );
  NAND2X1 U1835 ( .A(arr[895]), .B(n3428), .Y(n6466) );
  OAI21X1 U1836 ( .A(n5561), .B(n3423), .C(n6467), .Y(n9198) );
  NAND2X1 U1837 ( .A(arr[896]), .B(n3428), .Y(n6467) );
  OAI21X1 U1838 ( .A(n5563), .B(n3423), .C(n6468), .Y(n9199) );
  NAND2X1 U1839 ( .A(arr[897]), .B(n3428), .Y(n6468) );
  OAI21X1 U1840 ( .A(n5565), .B(n3423), .C(n6469), .Y(n9200) );
  NAND2X1 U1841 ( .A(arr[898]), .B(n3428), .Y(n6469) );
  OAI21X1 U1842 ( .A(n5567), .B(n3423), .C(n6470), .Y(n9201) );
  NAND2X1 U1843 ( .A(arr[899]), .B(n3428), .Y(n6470) );
  OAI21X1 U1844 ( .A(n5569), .B(n3423), .C(n6471), .Y(n9202) );
  NAND2X1 U1845 ( .A(arr[900]), .B(n3426), .Y(n6471) );
  OAI21X1 U1846 ( .A(n5571), .B(n3423), .C(n6472), .Y(n9203) );
  NAND2X1 U1847 ( .A(arr[901]), .B(n3426), .Y(n6472) );
  NAND2X1 U1848 ( .A(n6430), .B(n5617), .Y(n6431) );
  OAI21X1 U1849 ( .A(n5491), .B(n3417), .C(n6474), .Y(n9204) );
  NAND2X1 U1850 ( .A(arr[902]), .B(n3420), .Y(n6474) );
  OAI21X1 U1851 ( .A(n5493), .B(n3417), .C(n6475), .Y(n9205) );
  NAND2X1 U1852 ( .A(arr[903]), .B(n3420), .Y(n6475) );
  OAI21X1 U1853 ( .A(n5495), .B(n3417), .C(n6476), .Y(n9206) );
  NAND2X1 U1854 ( .A(arr[904]), .B(n3420), .Y(n6476) );
  OAI21X1 U1855 ( .A(n5497), .B(n3417), .C(n6477), .Y(n9207) );
  NAND2X1 U1856 ( .A(arr[905]), .B(n3420), .Y(n6477) );
  OAI21X1 U1857 ( .A(n5499), .B(n3417), .C(n6478), .Y(n9208) );
  NAND2X1 U1858 ( .A(arr[906]), .B(n3420), .Y(n6478) );
  OAI21X1 U1859 ( .A(n5501), .B(n3418), .C(n6479), .Y(n9209) );
  NAND2X1 U1860 ( .A(arr[907]), .B(n3420), .Y(n6479) );
  OAI21X1 U1861 ( .A(n5503), .B(n3418), .C(n6480), .Y(n9210) );
  NAND2X1 U1862 ( .A(arr[908]), .B(n3420), .Y(n6480) );
  OAI21X1 U1863 ( .A(n5505), .B(n3418), .C(n6481), .Y(n9211) );
  NAND2X1 U1864 ( .A(arr[909]), .B(n3420), .Y(n6481) );
  OAI21X1 U1865 ( .A(n5507), .B(n3417), .C(n6482), .Y(n9212) );
  NAND2X1 U1866 ( .A(arr[910]), .B(n3420), .Y(n6482) );
  OAI21X1 U1867 ( .A(n5509), .B(n3418), .C(n6483), .Y(n9213) );
  NAND2X1 U1868 ( .A(arr[911]), .B(n3420), .Y(n6483) );
  OAI21X1 U1869 ( .A(n5511), .B(n3419), .C(n6484), .Y(n9214) );
  NAND2X1 U1870 ( .A(arr[912]), .B(n3420), .Y(n6484) );
  OAI21X1 U1871 ( .A(n5513), .B(n3419), .C(n6485), .Y(n9215) );
  NAND2X1 U1872 ( .A(arr[913]), .B(n3420), .Y(n6485) );
  OAI21X1 U1873 ( .A(n5515), .B(n3419), .C(n6486), .Y(n9216) );
  NAND2X1 U1874 ( .A(arr[914]), .B(n3420), .Y(n6486) );
  OAI21X1 U1875 ( .A(n5517), .B(n3418), .C(n6487), .Y(n9217) );
  NAND2X1 U1876 ( .A(arr[915]), .B(n3421), .Y(n6487) );
  OAI21X1 U1877 ( .A(n5519), .B(n3420), .C(n6488), .Y(n9218) );
  NAND2X1 U1878 ( .A(arr[916]), .B(n3421), .Y(n6488) );
  OAI21X1 U1879 ( .A(n5521), .B(n3420), .C(n6489), .Y(n9219) );
  NAND2X1 U1880 ( .A(arr[917]), .B(n3421), .Y(n6489) );
  OAI21X1 U1881 ( .A(n5523), .B(n3419), .C(n6490), .Y(n9220) );
  NAND2X1 U1882 ( .A(arr[918]), .B(n3421), .Y(n6490) );
  OAI21X1 U1883 ( .A(n5525), .B(n3419), .C(n6491), .Y(n9221) );
  NAND2X1 U1884 ( .A(arr[919]), .B(n3421), .Y(n6491) );
  OAI21X1 U1885 ( .A(n5527), .B(n3419), .C(n6492), .Y(n9222) );
  NAND2X1 U1886 ( .A(arr[920]), .B(n3421), .Y(n6492) );
  OAI21X1 U1887 ( .A(n5529), .B(n3419), .C(n6493), .Y(n9223) );
  NAND2X1 U1888 ( .A(arr[921]), .B(n3421), .Y(n6493) );
  OAI21X1 U1889 ( .A(n5531), .B(n3419), .C(n6494), .Y(n9224) );
  NAND2X1 U1890 ( .A(arr[922]), .B(n3421), .Y(n6494) );
  OAI21X1 U1891 ( .A(n5533), .B(n3419), .C(n6495), .Y(n9225) );
  NAND2X1 U1892 ( .A(arr[923]), .B(n3421), .Y(n6495) );
  OAI21X1 U1893 ( .A(n5535), .B(n3419), .C(n6496), .Y(n9226) );
  NAND2X1 U1894 ( .A(arr[924]), .B(n3421), .Y(n6496) );
  OAI21X1 U1895 ( .A(n5537), .B(n3419), .C(n6497), .Y(n9227) );
  NAND2X1 U1896 ( .A(arr[925]), .B(n3421), .Y(n6497) );
  OAI21X1 U1897 ( .A(n5539), .B(n3419), .C(n6498), .Y(n9228) );
  NAND2X1 U1898 ( .A(arr[926]), .B(n3421), .Y(n6498) );
  OAI21X1 U1899 ( .A(n5541), .B(n3419), .C(n6499), .Y(n9229) );
  NAND2X1 U1900 ( .A(arr[927]), .B(n3421), .Y(n6499) );
  OAI21X1 U1901 ( .A(n5543), .B(n3418), .C(n6500), .Y(n9230) );
  NAND2X1 U1902 ( .A(arr[928]), .B(n3421), .Y(n6500) );
  OAI21X1 U1903 ( .A(n5545), .B(n3418), .C(n6501), .Y(n9231) );
  NAND2X1 U1904 ( .A(arr[929]), .B(n3421), .Y(n6501) );
  OAI21X1 U1905 ( .A(n5547), .B(n3418), .C(n6502), .Y(n9232) );
  NAND2X1 U1906 ( .A(arr[930]), .B(n3421), .Y(n6502) );
  OAI21X1 U1907 ( .A(n5549), .B(n3418), .C(n6503), .Y(n9233) );
  NAND2X1 U1908 ( .A(arr[931]), .B(n3421), .Y(n6503) );
  OAI21X1 U1909 ( .A(n5551), .B(n3418), .C(n6504), .Y(n9234) );
  NAND2X1 U1910 ( .A(arr[932]), .B(n3422), .Y(n6504) );
  OAI21X1 U1911 ( .A(n5553), .B(n3418), .C(n6505), .Y(n9235) );
  NAND2X1 U1912 ( .A(arr[933]), .B(n3422), .Y(n6505) );
  OAI21X1 U1913 ( .A(n5555), .B(n3418), .C(n6506), .Y(n9236) );
  NAND2X1 U1914 ( .A(arr[934]), .B(n3422), .Y(n6506) );
  OAI21X1 U1915 ( .A(n5557), .B(n3418), .C(n6507), .Y(n9237) );
  NAND2X1 U1916 ( .A(arr[935]), .B(n3422), .Y(n6507) );
  OAI21X1 U1917 ( .A(n5559), .B(n3417), .C(n6508), .Y(n9238) );
  NAND2X1 U1918 ( .A(arr[936]), .B(n3422), .Y(n6508) );
  OAI21X1 U1919 ( .A(n5561), .B(n3417), .C(n6509), .Y(n9239) );
  NAND2X1 U1920 ( .A(arr[937]), .B(n3422), .Y(n6509) );
  OAI21X1 U1921 ( .A(n5563), .B(n3417), .C(n6510), .Y(n9240) );
  NAND2X1 U1922 ( .A(arr[938]), .B(n3422), .Y(n6510) );
  OAI21X1 U1923 ( .A(n5565), .B(n3417), .C(n6511), .Y(n9241) );
  NAND2X1 U1924 ( .A(arr[939]), .B(n3422), .Y(n6511) );
  OAI21X1 U1925 ( .A(n5567), .B(n3417), .C(n6512), .Y(n9242) );
  NAND2X1 U1926 ( .A(arr[940]), .B(n3422), .Y(n6512) );
  OAI21X1 U1927 ( .A(n5569), .B(n3417), .C(n6513), .Y(n9243) );
  NAND2X1 U1928 ( .A(arr[941]), .B(n3420), .Y(n6513) );
  OAI21X1 U1929 ( .A(n5571), .B(n3417), .C(n6514), .Y(n9244) );
  NAND2X1 U1930 ( .A(arr[942]), .B(n3420), .Y(n6514) );
  NAND2X1 U1931 ( .A(n6430), .B(n5660), .Y(n6473) );
  OAI21X1 U1932 ( .A(n5491), .B(n3411), .C(n6516), .Y(n9245) );
  NAND2X1 U1933 ( .A(arr[943]), .B(n3414), .Y(n6516) );
  OAI21X1 U1934 ( .A(n5493), .B(n3411), .C(n6517), .Y(n9246) );
  NAND2X1 U1935 ( .A(arr[944]), .B(n3414), .Y(n6517) );
  OAI21X1 U1936 ( .A(n5495), .B(n3411), .C(n6518), .Y(n9247) );
  NAND2X1 U1937 ( .A(arr[945]), .B(n3414), .Y(n6518) );
  OAI21X1 U1938 ( .A(n5497), .B(n3411), .C(n6519), .Y(n9248) );
  NAND2X1 U1939 ( .A(arr[946]), .B(n3414), .Y(n6519) );
  OAI21X1 U1940 ( .A(n5499), .B(n3411), .C(n6520), .Y(n9249) );
  NAND2X1 U1941 ( .A(arr[947]), .B(n3414), .Y(n6520) );
  OAI21X1 U1942 ( .A(n5501), .B(n3412), .C(n6521), .Y(n9250) );
  NAND2X1 U1943 ( .A(arr[948]), .B(n3414), .Y(n6521) );
  OAI21X1 U1944 ( .A(n5503), .B(n3412), .C(n6522), .Y(n9251) );
  NAND2X1 U1945 ( .A(arr[949]), .B(n3414), .Y(n6522) );
  OAI21X1 U1946 ( .A(n5505), .B(n3412), .C(n6523), .Y(n9252) );
  NAND2X1 U1947 ( .A(arr[950]), .B(n3414), .Y(n6523) );
  OAI21X1 U1948 ( .A(n5507), .B(n3411), .C(n6524), .Y(n9253) );
  NAND2X1 U1949 ( .A(arr[951]), .B(n3414), .Y(n6524) );
  OAI21X1 U1950 ( .A(n5509), .B(n3412), .C(n6525), .Y(n9254) );
  NAND2X1 U1951 ( .A(arr[952]), .B(n3414), .Y(n6525) );
  OAI21X1 U1952 ( .A(n5511), .B(n3413), .C(n6526), .Y(n9255) );
  NAND2X1 U1953 ( .A(arr[953]), .B(n3414), .Y(n6526) );
  OAI21X1 U1954 ( .A(n5513), .B(n3413), .C(n6527), .Y(n9256) );
  NAND2X1 U1955 ( .A(arr[954]), .B(n3414), .Y(n6527) );
  OAI21X1 U1956 ( .A(n5515), .B(n3413), .C(n6528), .Y(n9257) );
  NAND2X1 U1957 ( .A(arr[955]), .B(n3414), .Y(n6528) );
  OAI21X1 U1958 ( .A(n5517), .B(n3412), .C(n6529), .Y(n9258) );
  NAND2X1 U1959 ( .A(arr[956]), .B(n3415), .Y(n6529) );
  OAI21X1 U1960 ( .A(n5519), .B(n3414), .C(n6530), .Y(n9259) );
  NAND2X1 U1961 ( .A(arr[957]), .B(n3415), .Y(n6530) );
  OAI21X1 U1962 ( .A(n5521), .B(n3414), .C(n6531), .Y(n9260) );
  NAND2X1 U1963 ( .A(arr[958]), .B(n3415), .Y(n6531) );
  OAI21X1 U1964 ( .A(n5523), .B(n3413), .C(n6532), .Y(n9261) );
  NAND2X1 U1965 ( .A(arr[959]), .B(n3415), .Y(n6532) );
  OAI21X1 U1966 ( .A(n5525), .B(n3413), .C(n6533), .Y(n9262) );
  NAND2X1 U1967 ( .A(arr[960]), .B(n3415), .Y(n6533) );
  OAI21X1 U1968 ( .A(n5527), .B(n3413), .C(n6534), .Y(n9263) );
  NAND2X1 U1969 ( .A(arr[961]), .B(n3415), .Y(n6534) );
  OAI21X1 U1970 ( .A(n5529), .B(n3413), .C(n6535), .Y(n9264) );
  NAND2X1 U1971 ( .A(arr[962]), .B(n3415), .Y(n6535) );
  OAI21X1 U1972 ( .A(n5531), .B(n3413), .C(n6536), .Y(n9265) );
  NAND2X1 U1973 ( .A(arr[963]), .B(n3415), .Y(n6536) );
  OAI21X1 U1974 ( .A(n5533), .B(n3413), .C(n6537), .Y(n9266) );
  NAND2X1 U1975 ( .A(arr[964]), .B(n3415), .Y(n6537) );
  OAI21X1 U1976 ( .A(n5535), .B(n3413), .C(n6538), .Y(n9267) );
  NAND2X1 U1977 ( .A(arr[965]), .B(n3415), .Y(n6538) );
  OAI21X1 U1978 ( .A(n5537), .B(n3413), .C(n6539), .Y(n9268) );
  NAND2X1 U1979 ( .A(arr[966]), .B(n3415), .Y(n6539) );
  OAI21X1 U1980 ( .A(n5539), .B(n3413), .C(n6540), .Y(n9269) );
  NAND2X1 U1981 ( .A(arr[967]), .B(n3415), .Y(n6540) );
  OAI21X1 U1982 ( .A(n5541), .B(n3413), .C(n6541), .Y(n9270) );
  NAND2X1 U1983 ( .A(arr[968]), .B(n3415), .Y(n6541) );
  OAI21X1 U1984 ( .A(n5543), .B(n3412), .C(n6542), .Y(n9271) );
  NAND2X1 U1985 ( .A(arr[969]), .B(n3415), .Y(n6542) );
  OAI21X1 U1986 ( .A(n5545), .B(n3412), .C(n6543), .Y(n9272) );
  NAND2X1 U1987 ( .A(arr[970]), .B(n3415), .Y(n6543) );
  OAI21X1 U1988 ( .A(n5547), .B(n3412), .C(n6544), .Y(n9273) );
  NAND2X1 U1989 ( .A(arr[971]), .B(n3415), .Y(n6544) );
  OAI21X1 U1990 ( .A(n5549), .B(n3412), .C(n6545), .Y(n9274) );
  NAND2X1 U1991 ( .A(arr[972]), .B(n3415), .Y(n6545) );
  OAI21X1 U1992 ( .A(n5551), .B(n3412), .C(n6546), .Y(n9275) );
  NAND2X1 U1993 ( .A(arr[973]), .B(n3416), .Y(n6546) );
  OAI21X1 U1994 ( .A(n5553), .B(n3412), .C(n6547), .Y(n9276) );
  NAND2X1 U1995 ( .A(arr[974]), .B(n3416), .Y(n6547) );
  OAI21X1 U1996 ( .A(n5555), .B(n3412), .C(n6548), .Y(n9277) );
  NAND2X1 U1997 ( .A(arr[975]), .B(n3416), .Y(n6548) );
  OAI21X1 U1998 ( .A(n5557), .B(n3412), .C(n6549), .Y(n9278) );
  NAND2X1 U1999 ( .A(arr[976]), .B(n3416), .Y(n6549) );
  OAI21X1 U2000 ( .A(n5559), .B(n3411), .C(n6550), .Y(n9279) );
  NAND2X1 U2001 ( .A(arr[977]), .B(n3416), .Y(n6550) );
  OAI21X1 U2002 ( .A(n5561), .B(n3411), .C(n6551), .Y(n9280) );
  NAND2X1 U2003 ( .A(arr[978]), .B(n3416), .Y(n6551) );
  OAI21X1 U2004 ( .A(n5563), .B(n3411), .C(n6552), .Y(n9281) );
  NAND2X1 U2005 ( .A(arr[979]), .B(n3416), .Y(n6552) );
  OAI21X1 U2006 ( .A(n5565), .B(n3411), .C(n6553), .Y(n9282) );
  NAND2X1 U2007 ( .A(arr[980]), .B(n3416), .Y(n6553) );
  OAI21X1 U2008 ( .A(n5567), .B(n3411), .C(n6554), .Y(n9283) );
  NAND2X1 U2009 ( .A(arr[981]), .B(n3416), .Y(n6554) );
  OAI21X1 U2010 ( .A(n5569), .B(n3411), .C(n6555), .Y(n9284) );
  NAND2X1 U2011 ( .A(arr[982]), .B(n3414), .Y(n6555) );
  OAI21X1 U2012 ( .A(n5571), .B(n3411), .C(n6556), .Y(n9285) );
  NAND2X1 U2013 ( .A(arr[983]), .B(n3414), .Y(n6556) );
  NAND2X1 U2014 ( .A(n6430), .B(n5703), .Y(n6515) );
  OAI21X1 U2016 ( .A(n5491), .B(n3405), .C(n6558), .Y(n9286) );
  NAND2X1 U2017 ( .A(arr[984]), .B(n3408), .Y(n6558) );
  OAI21X1 U2018 ( .A(n5493), .B(n3405), .C(n6559), .Y(n9287) );
  NAND2X1 U2019 ( .A(arr[985]), .B(n3408), .Y(n6559) );
  OAI21X1 U2020 ( .A(n5495), .B(n3405), .C(n6560), .Y(n9288) );
  NAND2X1 U2021 ( .A(arr[986]), .B(n3408), .Y(n6560) );
  OAI21X1 U2022 ( .A(n5497), .B(n3405), .C(n6561), .Y(n9289) );
  NAND2X1 U2023 ( .A(arr[987]), .B(n3408), .Y(n6561) );
  OAI21X1 U2024 ( .A(n5499), .B(n3405), .C(n6562), .Y(n9290) );
  NAND2X1 U2025 ( .A(arr[988]), .B(n3408), .Y(n6562) );
  OAI21X1 U2026 ( .A(n5501), .B(n3406), .C(n6563), .Y(n9291) );
  NAND2X1 U2027 ( .A(arr[989]), .B(n3408), .Y(n6563) );
  OAI21X1 U2028 ( .A(n5503), .B(n3406), .C(n6564), .Y(n9292) );
  NAND2X1 U2029 ( .A(arr[990]), .B(n3408), .Y(n6564) );
  OAI21X1 U2030 ( .A(n5505), .B(n3406), .C(n6565), .Y(n9293) );
  NAND2X1 U2031 ( .A(arr[991]), .B(n3408), .Y(n6565) );
  OAI21X1 U2032 ( .A(n5507), .B(n3405), .C(n6566), .Y(n9294) );
  NAND2X1 U2033 ( .A(arr[992]), .B(n3408), .Y(n6566) );
  OAI21X1 U2034 ( .A(n5509), .B(n3406), .C(n6567), .Y(n9295) );
  NAND2X1 U2035 ( .A(arr[993]), .B(n3408), .Y(n6567) );
  OAI21X1 U2036 ( .A(n5511), .B(n3407), .C(n6568), .Y(n9296) );
  NAND2X1 U2037 ( .A(arr[994]), .B(n3408), .Y(n6568) );
  OAI21X1 U2038 ( .A(n5513), .B(n3407), .C(n6569), .Y(n9297) );
  NAND2X1 U2039 ( .A(arr[995]), .B(n3408), .Y(n6569) );
  OAI21X1 U2040 ( .A(n5515), .B(n3407), .C(n6570), .Y(n9298) );
  NAND2X1 U2041 ( .A(arr[996]), .B(n3408), .Y(n6570) );
  OAI21X1 U2042 ( .A(n5517), .B(n3406), .C(n6571), .Y(n9299) );
  NAND2X1 U2043 ( .A(arr[997]), .B(n3409), .Y(n6571) );
  OAI21X1 U2044 ( .A(n5519), .B(n3408), .C(n6572), .Y(n9300) );
  NAND2X1 U2045 ( .A(arr[998]), .B(n3409), .Y(n6572) );
  OAI21X1 U2046 ( .A(n5521), .B(n3408), .C(n6573), .Y(n9301) );
  NAND2X1 U2047 ( .A(arr[999]), .B(n3409), .Y(n6573) );
  OAI21X1 U2048 ( .A(n5523), .B(n3407), .C(n6574), .Y(n9302) );
  NAND2X1 U2049 ( .A(arr[1000]), .B(n3409), .Y(n6574) );
  OAI21X1 U2050 ( .A(n5525), .B(n3407), .C(n6575), .Y(n9303) );
  NAND2X1 U2051 ( .A(arr[1001]), .B(n3409), .Y(n6575) );
  OAI21X1 U2052 ( .A(n5527), .B(n3407), .C(n6576), .Y(n9304) );
  NAND2X1 U2053 ( .A(arr[1002]), .B(n3409), .Y(n6576) );
  OAI21X1 U2054 ( .A(n5529), .B(n3407), .C(n6577), .Y(n9305) );
  NAND2X1 U2055 ( .A(arr[1003]), .B(n3409), .Y(n6577) );
  OAI21X1 U2056 ( .A(n5531), .B(n3407), .C(n6578), .Y(n9306) );
  NAND2X1 U2057 ( .A(arr[1004]), .B(n3409), .Y(n6578) );
  OAI21X1 U2058 ( .A(n5533), .B(n3407), .C(n6579), .Y(n9307) );
  NAND2X1 U2059 ( .A(arr[1005]), .B(n3409), .Y(n6579) );
  OAI21X1 U2060 ( .A(n5535), .B(n3407), .C(n6580), .Y(n9308) );
  NAND2X1 U2061 ( .A(arr[1006]), .B(n3409), .Y(n6580) );
  OAI21X1 U2062 ( .A(n5537), .B(n3407), .C(n6581), .Y(n9309) );
  NAND2X1 U2063 ( .A(arr[1007]), .B(n3409), .Y(n6581) );
  OAI21X1 U2064 ( .A(n5539), .B(n3407), .C(n6582), .Y(n9310) );
  NAND2X1 U2065 ( .A(arr[1008]), .B(n3409), .Y(n6582) );
  OAI21X1 U2066 ( .A(n5541), .B(n3407), .C(n6583), .Y(n9311) );
  NAND2X1 U2067 ( .A(arr[1009]), .B(n3409), .Y(n6583) );
  OAI21X1 U2068 ( .A(n5543), .B(n3406), .C(n6584), .Y(n9312) );
  NAND2X1 U2069 ( .A(arr[1010]), .B(n3409), .Y(n6584) );
  OAI21X1 U2070 ( .A(n5545), .B(n3406), .C(n6585), .Y(n9313) );
  NAND2X1 U2071 ( .A(arr[1011]), .B(n3409), .Y(n6585) );
  OAI21X1 U2072 ( .A(n5547), .B(n3406), .C(n6586), .Y(n9314) );
  NAND2X1 U2073 ( .A(arr[1012]), .B(n3409), .Y(n6586) );
  OAI21X1 U2074 ( .A(n5549), .B(n3406), .C(n6587), .Y(n9315) );
  NAND2X1 U2075 ( .A(arr[1013]), .B(n3409), .Y(n6587) );
  OAI21X1 U2076 ( .A(n5551), .B(n3406), .C(n6588), .Y(n9316) );
  NAND2X1 U2077 ( .A(arr[1014]), .B(n3410), .Y(n6588) );
  OAI21X1 U2078 ( .A(n5553), .B(n3406), .C(n6589), .Y(n9317) );
  NAND2X1 U2079 ( .A(arr[1015]), .B(n3410), .Y(n6589) );
  OAI21X1 U2080 ( .A(n5555), .B(n3406), .C(n6590), .Y(n9318) );
  NAND2X1 U2081 ( .A(arr[1016]), .B(n3410), .Y(n6590) );
  OAI21X1 U2082 ( .A(n5557), .B(n3406), .C(n6591), .Y(n9319) );
  NAND2X1 U2083 ( .A(arr[1017]), .B(n3410), .Y(n6591) );
  OAI21X1 U2084 ( .A(n5559), .B(n3405), .C(n6592), .Y(n9320) );
  NAND2X1 U2085 ( .A(arr[1018]), .B(n3410), .Y(n6592) );
  OAI21X1 U2086 ( .A(n5561), .B(n3405), .C(n6593), .Y(n9321) );
  NAND2X1 U2087 ( .A(arr[1019]), .B(n3410), .Y(n6593) );
  OAI21X1 U2088 ( .A(n5563), .B(n3405), .C(n6594), .Y(n9322) );
  NAND2X1 U2089 ( .A(arr[1020]), .B(n3410), .Y(n6594) );
  OAI21X1 U2090 ( .A(n5565), .B(n3405), .C(n6595), .Y(n9323) );
  NAND2X1 U2091 ( .A(arr[1021]), .B(n3410), .Y(n6595) );
  OAI21X1 U2092 ( .A(n5567), .B(n3405), .C(n6596), .Y(n9324) );
  NAND2X1 U2093 ( .A(arr[1022]), .B(n3410), .Y(n6596) );
  OAI21X1 U2094 ( .A(n5569), .B(n3405), .C(n6597), .Y(n9325) );
  NAND2X1 U2095 ( .A(arr[1023]), .B(n3408), .Y(n6597) );
  OAI21X1 U2096 ( .A(n5571), .B(n3405), .C(n6598), .Y(n9326) );
  NAND2X1 U2097 ( .A(arr[1024]), .B(n3408), .Y(n6598) );
  NAND2X1 U2098 ( .A(n6599), .B(n5573), .Y(n6557) );
  OAI21X1 U2099 ( .A(n5491), .B(n3399), .C(n6601), .Y(n9327) );
  NAND2X1 U2100 ( .A(arr[1025]), .B(n3402), .Y(n6601) );
  OAI21X1 U2101 ( .A(n5493), .B(n3399), .C(n6602), .Y(n9328) );
  NAND2X1 U2102 ( .A(arr[1026]), .B(n3402), .Y(n6602) );
  OAI21X1 U2103 ( .A(n5495), .B(n3399), .C(n6603), .Y(n9329) );
  NAND2X1 U2104 ( .A(arr[1027]), .B(n3402), .Y(n6603) );
  OAI21X1 U2105 ( .A(n5497), .B(n3399), .C(n6604), .Y(n9330) );
  NAND2X1 U2106 ( .A(arr[1028]), .B(n3402), .Y(n6604) );
  OAI21X1 U2107 ( .A(n5499), .B(n3399), .C(n6605), .Y(n9331) );
  NAND2X1 U2108 ( .A(arr[1029]), .B(n3402), .Y(n6605) );
  OAI21X1 U2109 ( .A(n5501), .B(n3400), .C(n6606), .Y(n9332) );
  NAND2X1 U2110 ( .A(arr[1030]), .B(n3402), .Y(n6606) );
  OAI21X1 U2111 ( .A(n5503), .B(n3400), .C(n6607), .Y(n9333) );
  NAND2X1 U2112 ( .A(arr[1031]), .B(n3402), .Y(n6607) );
  OAI21X1 U2113 ( .A(n5505), .B(n3400), .C(n6608), .Y(n9334) );
  NAND2X1 U2114 ( .A(arr[1032]), .B(n3402), .Y(n6608) );
  OAI21X1 U2115 ( .A(n5507), .B(n3399), .C(n6609), .Y(n9335) );
  NAND2X1 U2116 ( .A(arr[1033]), .B(n3402), .Y(n6609) );
  OAI21X1 U2117 ( .A(n5509), .B(n3400), .C(n6610), .Y(n9336) );
  NAND2X1 U2118 ( .A(arr[1034]), .B(n3402), .Y(n6610) );
  OAI21X1 U2119 ( .A(n5511), .B(n3401), .C(n6611), .Y(n9337) );
  NAND2X1 U2120 ( .A(arr[1035]), .B(n3402), .Y(n6611) );
  OAI21X1 U2121 ( .A(n5513), .B(n3401), .C(n6612), .Y(n9338) );
  NAND2X1 U2122 ( .A(arr[1036]), .B(n3402), .Y(n6612) );
  OAI21X1 U2123 ( .A(n5515), .B(n3401), .C(n6613), .Y(n9339) );
  NAND2X1 U2124 ( .A(arr[1037]), .B(n3402), .Y(n6613) );
  OAI21X1 U2125 ( .A(n5517), .B(n3400), .C(n6614), .Y(n9340) );
  NAND2X1 U2126 ( .A(arr[1038]), .B(n3403), .Y(n6614) );
  OAI21X1 U2127 ( .A(n5519), .B(n3402), .C(n6615), .Y(n9341) );
  NAND2X1 U2128 ( .A(arr[1039]), .B(n3403), .Y(n6615) );
  OAI21X1 U2129 ( .A(n5521), .B(n3402), .C(n6616), .Y(n9342) );
  NAND2X1 U2130 ( .A(arr[1040]), .B(n3403), .Y(n6616) );
  OAI21X1 U2131 ( .A(n5523), .B(n3401), .C(n6617), .Y(n9343) );
  NAND2X1 U2132 ( .A(arr[1041]), .B(n3403), .Y(n6617) );
  OAI21X1 U2133 ( .A(n5525), .B(n3401), .C(n6618), .Y(n9344) );
  NAND2X1 U2134 ( .A(arr[1042]), .B(n3403), .Y(n6618) );
  OAI21X1 U2135 ( .A(n5527), .B(n3401), .C(n6619), .Y(n9345) );
  NAND2X1 U2136 ( .A(arr[1043]), .B(n3403), .Y(n6619) );
  OAI21X1 U2137 ( .A(n5529), .B(n3401), .C(n6620), .Y(n9346) );
  NAND2X1 U2138 ( .A(arr[1044]), .B(n3403), .Y(n6620) );
  OAI21X1 U2139 ( .A(n5531), .B(n3401), .C(n6621), .Y(n9347) );
  NAND2X1 U2140 ( .A(arr[1045]), .B(n3403), .Y(n6621) );
  OAI21X1 U2141 ( .A(n5533), .B(n3401), .C(n6622), .Y(n9348) );
  NAND2X1 U2142 ( .A(arr[1046]), .B(n3403), .Y(n6622) );
  OAI21X1 U2143 ( .A(n5535), .B(n3401), .C(n6623), .Y(n9349) );
  NAND2X1 U2144 ( .A(arr[1047]), .B(n3403), .Y(n6623) );
  OAI21X1 U2145 ( .A(n5537), .B(n3401), .C(n6624), .Y(n9350) );
  NAND2X1 U2146 ( .A(arr[1048]), .B(n3403), .Y(n6624) );
  OAI21X1 U2147 ( .A(n5539), .B(n3401), .C(n6625), .Y(n9351) );
  NAND2X1 U2148 ( .A(arr[1049]), .B(n3403), .Y(n6625) );
  OAI21X1 U2149 ( .A(n5541), .B(n3401), .C(n6626), .Y(n9352) );
  NAND2X1 U2150 ( .A(arr[1050]), .B(n3403), .Y(n6626) );
  OAI21X1 U2151 ( .A(n5543), .B(n3400), .C(n6627), .Y(n9353) );
  NAND2X1 U2152 ( .A(arr[1051]), .B(n3403), .Y(n6627) );
  OAI21X1 U2153 ( .A(n5545), .B(n3400), .C(n6628), .Y(n9354) );
  NAND2X1 U2154 ( .A(arr[1052]), .B(n3403), .Y(n6628) );
  OAI21X1 U2155 ( .A(n5547), .B(n3400), .C(n6629), .Y(n9355) );
  NAND2X1 U2156 ( .A(arr[1053]), .B(n3403), .Y(n6629) );
  OAI21X1 U2157 ( .A(n5549), .B(n3400), .C(n6630), .Y(n9356) );
  NAND2X1 U2158 ( .A(arr[1054]), .B(n3403), .Y(n6630) );
  OAI21X1 U2159 ( .A(n5551), .B(n3400), .C(n6631), .Y(n9357) );
  NAND2X1 U2160 ( .A(arr[1055]), .B(n3404), .Y(n6631) );
  OAI21X1 U2161 ( .A(n5553), .B(n3400), .C(n6632), .Y(n9358) );
  NAND2X1 U2162 ( .A(arr[1056]), .B(n3404), .Y(n6632) );
  OAI21X1 U2163 ( .A(n5555), .B(n3400), .C(n6633), .Y(n9359) );
  NAND2X1 U2164 ( .A(arr[1057]), .B(n3404), .Y(n6633) );
  OAI21X1 U2165 ( .A(n5557), .B(n3400), .C(n6634), .Y(n9360) );
  NAND2X1 U2166 ( .A(arr[1058]), .B(n3404), .Y(n6634) );
  OAI21X1 U2167 ( .A(n5559), .B(n3399), .C(n6635), .Y(n9361) );
  NAND2X1 U2168 ( .A(arr[1059]), .B(n3404), .Y(n6635) );
  OAI21X1 U2169 ( .A(n5561), .B(n3399), .C(n6636), .Y(n9362) );
  NAND2X1 U2170 ( .A(arr[1060]), .B(n3404), .Y(n6636) );
  OAI21X1 U2171 ( .A(n5563), .B(n3399), .C(n6637), .Y(n9363) );
  NAND2X1 U2172 ( .A(arr[1061]), .B(n3404), .Y(n6637) );
  OAI21X1 U2173 ( .A(n5565), .B(n3399), .C(n6638), .Y(n9364) );
  NAND2X1 U2174 ( .A(arr[1062]), .B(n3404), .Y(n6638) );
  OAI21X1 U2175 ( .A(n5567), .B(n3399), .C(n6639), .Y(n9365) );
  NAND2X1 U2176 ( .A(arr[1063]), .B(n3404), .Y(n6639) );
  OAI21X1 U2177 ( .A(n5569), .B(n3399), .C(n6640), .Y(n9366) );
  NAND2X1 U2178 ( .A(arr[1064]), .B(n3402), .Y(n6640) );
  OAI21X1 U2179 ( .A(n5571), .B(n3399), .C(n6641), .Y(n9367) );
  NAND2X1 U2180 ( .A(arr[1065]), .B(n3402), .Y(n6641) );
  NAND2X1 U2181 ( .A(n6599), .B(n5617), .Y(n6600) );
  OAI21X1 U2182 ( .A(n5491), .B(n3393), .C(n6643), .Y(n9368) );
  NAND2X1 U2183 ( .A(arr[1066]), .B(n3396), .Y(n6643) );
  OAI21X1 U2184 ( .A(n5493), .B(n3393), .C(n6644), .Y(n9369) );
  NAND2X1 U2185 ( .A(arr[1067]), .B(n3396), .Y(n6644) );
  OAI21X1 U2186 ( .A(n5495), .B(n3393), .C(n6645), .Y(n9370) );
  NAND2X1 U2187 ( .A(arr[1068]), .B(n3396), .Y(n6645) );
  OAI21X1 U2188 ( .A(n5497), .B(n3393), .C(n6646), .Y(n9371) );
  NAND2X1 U2189 ( .A(arr[1069]), .B(n3396), .Y(n6646) );
  OAI21X1 U2190 ( .A(n5499), .B(n3393), .C(n6647), .Y(n9372) );
  NAND2X1 U2191 ( .A(arr[1070]), .B(n3396), .Y(n6647) );
  OAI21X1 U2192 ( .A(n5501), .B(n3394), .C(n6648), .Y(n9373) );
  NAND2X1 U2193 ( .A(arr[1071]), .B(n3396), .Y(n6648) );
  OAI21X1 U2194 ( .A(n5503), .B(n3394), .C(n6649), .Y(n9374) );
  NAND2X1 U2195 ( .A(arr[1072]), .B(n3396), .Y(n6649) );
  OAI21X1 U2196 ( .A(n5505), .B(n3394), .C(n6650), .Y(n9375) );
  NAND2X1 U2197 ( .A(arr[1073]), .B(n3396), .Y(n6650) );
  OAI21X1 U2198 ( .A(n5507), .B(n3393), .C(n6651), .Y(n9376) );
  NAND2X1 U2199 ( .A(arr[1074]), .B(n3396), .Y(n6651) );
  OAI21X1 U2200 ( .A(n5509), .B(n3394), .C(n6652), .Y(n9377) );
  NAND2X1 U2201 ( .A(arr[1075]), .B(n3396), .Y(n6652) );
  OAI21X1 U2202 ( .A(n5511), .B(n3395), .C(n6653), .Y(n9378) );
  NAND2X1 U2203 ( .A(arr[1076]), .B(n3396), .Y(n6653) );
  OAI21X1 U2204 ( .A(n5513), .B(n3395), .C(n6654), .Y(n9379) );
  NAND2X1 U2205 ( .A(arr[1077]), .B(n3396), .Y(n6654) );
  OAI21X1 U2206 ( .A(n5515), .B(n3395), .C(n6655), .Y(n9380) );
  NAND2X1 U2207 ( .A(arr[1078]), .B(n3396), .Y(n6655) );
  OAI21X1 U2208 ( .A(n5517), .B(n3394), .C(n6656), .Y(n9381) );
  NAND2X1 U2209 ( .A(arr[1079]), .B(n3397), .Y(n6656) );
  OAI21X1 U2210 ( .A(n5519), .B(n3396), .C(n6657), .Y(n9382) );
  NAND2X1 U2211 ( .A(arr[1080]), .B(n3397), .Y(n6657) );
  OAI21X1 U2212 ( .A(n5521), .B(n3396), .C(n6658), .Y(n9383) );
  NAND2X1 U2213 ( .A(arr[1081]), .B(n3397), .Y(n6658) );
  OAI21X1 U2214 ( .A(n5523), .B(n3395), .C(n6659), .Y(n9384) );
  NAND2X1 U2215 ( .A(arr[1082]), .B(n3397), .Y(n6659) );
  OAI21X1 U2216 ( .A(n5525), .B(n3395), .C(n6660), .Y(n9385) );
  NAND2X1 U2217 ( .A(arr[1083]), .B(n3397), .Y(n6660) );
  OAI21X1 U2218 ( .A(n5527), .B(n3395), .C(n6661), .Y(n9386) );
  NAND2X1 U2219 ( .A(arr[1084]), .B(n3397), .Y(n6661) );
  OAI21X1 U2220 ( .A(n5529), .B(n3395), .C(n6662), .Y(n9387) );
  NAND2X1 U2221 ( .A(arr[1085]), .B(n3397), .Y(n6662) );
  OAI21X1 U2222 ( .A(n5531), .B(n3395), .C(n6663), .Y(n9388) );
  NAND2X1 U2223 ( .A(arr[1086]), .B(n3397), .Y(n6663) );
  OAI21X1 U2224 ( .A(n5533), .B(n3395), .C(n6664), .Y(n9389) );
  NAND2X1 U2225 ( .A(arr[1087]), .B(n3397), .Y(n6664) );
  OAI21X1 U2226 ( .A(n5535), .B(n3395), .C(n6665), .Y(n9390) );
  NAND2X1 U2227 ( .A(arr[1088]), .B(n3397), .Y(n6665) );
  OAI21X1 U2228 ( .A(n5537), .B(n3395), .C(n6666), .Y(n9391) );
  NAND2X1 U2229 ( .A(arr[1089]), .B(n3397), .Y(n6666) );
  OAI21X1 U2230 ( .A(n5539), .B(n3395), .C(n6667), .Y(n9392) );
  NAND2X1 U2231 ( .A(arr[1090]), .B(n3397), .Y(n6667) );
  OAI21X1 U2232 ( .A(n5541), .B(n3395), .C(n6668), .Y(n9393) );
  NAND2X1 U2233 ( .A(arr[1091]), .B(n3397), .Y(n6668) );
  OAI21X1 U2234 ( .A(n5543), .B(n3394), .C(n6669), .Y(n9394) );
  NAND2X1 U2235 ( .A(arr[1092]), .B(n3397), .Y(n6669) );
  OAI21X1 U2236 ( .A(n5545), .B(n3394), .C(n6670), .Y(n9395) );
  NAND2X1 U2237 ( .A(arr[1093]), .B(n3397), .Y(n6670) );
  OAI21X1 U2238 ( .A(n5547), .B(n3394), .C(n6671), .Y(n9396) );
  NAND2X1 U2239 ( .A(arr[1094]), .B(n3397), .Y(n6671) );
  OAI21X1 U2240 ( .A(n5549), .B(n3394), .C(n6672), .Y(n9397) );
  NAND2X1 U2241 ( .A(arr[1095]), .B(n3397), .Y(n6672) );
  OAI21X1 U2242 ( .A(n5551), .B(n3394), .C(n6673), .Y(n9398) );
  NAND2X1 U2243 ( .A(arr[1096]), .B(n3398), .Y(n6673) );
  OAI21X1 U2244 ( .A(n5553), .B(n3394), .C(n6674), .Y(n9399) );
  NAND2X1 U2245 ( .A(arr[1097]), .B(n3398), .Y(n6674) );
  OAI21X1 U2246 ( .A(n5555), .B(n3394), .C(n6675), .Y(n9400) );
  NAND2X1 U2247 ( .A(arr[1098]), .B(n3398), .Y(n6675) );
  OAI21X1 U2248 ( .A(n5557), .B(n3394), .C(n6676), .Y(n9401) );
  NAND2X1 U2249 ( .A(arr[1099]), .B(n3398), .Y(n6676) );
  OAI21X1 U2250 ( .A(n5559), .B(n3393), .C(n6677), .Y(n9402) );
  NAND2X1 U2251 ( .A(arr[1100]), .B(n3398), .Y(n6677) );
  OAI21X1 U2252 ( .A(n5561), .B(n3393), .C(n6678), .Y(n9403) );
  NAND2X1 U2253 ( .A(arr[1101]), .B(n3398), .Y(n6678) );
  OAI21X1 U2254 ( .A(n5563), .B(n3393), .C(n6679), .Y(n9404) );
  NAND2X1 U2255 ( .A(arr[1102]), .B(n3398), .Y(n6679) );
  OAI21X1 U2256 ( .A(n5565), .B(n3393), .C(n6680), .Y(n9405) );
  NAND2X1 U2257 ( .A(arr[1103]), .B(n3398), .Y(n6680) );
  OAI21X1 U2258 ( .A(n5567), .B(n3393), .C(n6681), .Y(n9406) );
  NAND2X1 U2259 ( .A(arr[1104]), .B(n3398), .Y(n6681) );
  OAI21X1 U2260 ( .A(n5569), .B(n3393), .C(n6682), .Y(n9407) );
  NAND2X1 U2261 ( .A(arr[1105]), .B(n3396), .Y(n6682) );
  OAI21X1 U2262 ( .A(n5571), .B(n3393), .C(n6683), .Y(n9408) );
  NAND2X1 U2263 ( .A(arr[1106]), .B(n3396), .Y(n6683) );
  NAND2X1 U2264 ( .A(n6599), .B(n5660), .Y(n6642) );
  OAI21X1 U2265 ( .A(n5491), .B(n3387), .C(n6685), .Y(n9409) );
  NAND2X1 U2266 ( .A(arr[1107]), .B(n3390), .Y(n6685) );
  OAI21X1 U2267 ( .A(n5493), .B(n3387), .C(n6686), .Y(n9410) );
  NAND2X1 U2268 ( .A(arr[1108]), .B(n3390), .Y(n6686) );
  OAI21X1 U2269 ( .A(n5495), .B(n3387), .C(n6687), .Y(n9411) );
  NAND2X1 U2270 ( .A(arr[1109]), .B(n3390), .Y(n6687) );
  OAI21X1 U2271 ( .A(n5497), .B(n3387), .C(n6688), .Y(n9412) );
  NAND2X1 U2272 ( .A(arr[1110]), .B(n3390), .Y(n6688) );
  OAI21X1 U2273 ( .A(n5499), .B(n3387), .C(n6689), .Y(n9413) );
  NAND2X1 U2274 ( .A(arr[1111]), .B(n3390), .Y(n6689) );
  OAI21X1 U2275 ( .A(n5501), .B(n3388), .C(n6690), .Y(n9414) );
  NAND2X1 U2276 ( .A(arr[1112]), .B(n3390), .Y(n6690) );
  OAI21X1 U2277 ( .A(n5503), .B(n3388), .C(n6691), .Y(n9415) );
  NAND2X1 U2278 ( .A(arr[1113]), .B(n3390), .Y(n6691) );
  OAI21X1 U2279 ( .A(n5505), .B(n3388), .C(n6692), .Y(n9416) );
  NAND2X1 U2280 ( .A(arr[1114]), .B(n3390), .Y(n6692) );
  OAI21X1 U2281 ( .A(n5507), .B(n3387), .C(n6693), .Y(n9417) );
  NAND2X1 U2282 ( .A(arr[1115]), .B(n3390), .Y(n6693) );
  OAI21X1 U2283 ( .A(n5509), .B(n3388), .C(n6694), .Y(n9418) );
  NAND2X1 U2284 ( .A(arr[1116]), .B(n3390), .Y(n6694) );
  OAI21X1 U2285 ( .A(n5511), .B(n3389), .C(n6695), .Y(n9419) );
  NAND2X1 U2286 ( .A(arr[1117]), .B(n3390), .Y(n6695) );
  OAI21X1 U2287 ( .A(n5513), .B(n3389), .C(n6696), .Y(n9420) );
  NAND2X1 U2288 ( .A(arr[1118]), .B(n3390), .Y(n6696) );
  OAI21X1 U2289 ( .A(n5515), .B(n3389), .C(n6697), .Y(n9421) );
  NAND2X1 U2290 ( .A(arr[1119]), .B(n3390), .Y(n6697) );
  OAI21X1 U2291 ( .A(n5517), .B(n3388), .C(n6698), .Y(n9422) );
  NAND2X1 U2292 ( .A(arr[1120]), .B(n3391), .Y(n6698) );
  OAI21X1 U2293 ( .A(n5519), .B(n3390), .C(n6699), .Y(n9423) );
  NAND2X1 U2294 ( .A(arr[1121]), .B(n3391), .Y(n6699) );
  OAI21X1 U2295 ( .A(n5521), .B(n3390), .C(n6700), .Y(n9424) );
  NAND2X1 U2296 ( .A(arr[1122]), .B(n3391), .Y(n6700) );
  OAI21X1 U2297 ( .A(n5523), .B(n3389), .C(n6701), .Y(n9425) );
  NAND2X1 U2298 ( .A(arr[1123]), .B(n3391), .Y(n6701) );
  OAI21X1 U2299 ( .A(n5525), .B(n3389), .C(n6702), .Y(n9426) );
  NAND2X1 U2300 ( .A(arr[1124]), .B(n3391), .Y(n6702) );
  OAI21X1 U2301 ( .A(n5527), .B(n3389), .C(n6703), .Y(n9427) );
  NAND2X1 U2302 ( .A(arr[1125]), .B(n3391), .Y(n6703) );
  OAI21X1 U2303 ( .A(n5529), .B(n3389), .C(n6704), .Y(n9428) );
  NAND2X1 U2304 ( .A(arr[1126]), .B(n3391), .Y(n6704) );
  OAI21X1 U2305 ( .A(n5531), .B(n3389), .C(n6705), .Y(n9429) );
  NAND2X1 U2306 ( .A(arr[1127]), .B(n3391), .Y(n6705) );
  OAI21X1 U2307 ( .A(n5533), .B(n3389), .C(n6706), .Y(n9430) );
  NAND2X1 U2308 ( .A(arr[1128]), .B(n3391), .Y(n6706) );
  OAI21X1 U2309 ( .A(n5535), .B(n3389), .C(n6707), .Y(n9431) );
  NAND2X1 U2310 ( .A(arr[1129]), .B(n3391), .Y(n6707) );
  OAI21X1 U2311 ( .A(n5537), .B(n3389), .C(n6708), .Y(n9432) );
  NAND2X1 U2312 ( .A(arr[1130]), .B(n3391), .Y(n6708) );
  OAI21X1 U2313 ( .A(n5539), .B(n3389), .C(n6709), .Y(n9433) );
  NAND2X1 U2314 ( .A(arr[1131]), .B(n3391), .Y(n6709) );
  OAI21X1 U2315 ( .A(n5541), .B(n3389), .C(n6710), .Y(n9434) );
  NAND2X1 U2316 ( .A(arr[1132]), .B(n3391), .Y(n6710) );
  OAI21X1 U2317 ( .A(n5543), .B(n3388), .C(n6711), .Y(n9435) );
  NAND2X1 U2318 ( .A(arr[1133]), .B(n3391), .Y(n6711) );
  OAI21X1 U2319 ( .A(n5545), .B(n3388), .C(n6712), .Y(n9436) );
  NAND2X1 U2320 ( .A(arr[1134]), .B(n3391), .Y(n6712) );
  OAI21X1 U2321 ( .A(n5547), .B(n3388), .C(n6713), .Y(n9437) );
  NAND2X1 U2322 ( .A(arr[1135]), .B(n3391), .Y(n6713) );
  OAI21X1 U2323 ( .A(n5549), .B(n3388), .C(n6714), .Y(n9438) );
  NAND2X1 U2324 ( .A(arr[1136]), .B(n3391), .Y(n6714) );
  OAI21X1 U2325 ( .A(n5551), .B(n3388), .C(n6715), .Y(n9439) );
  NAND2X1 U2326 ( .A(arr[1137]), .B(n3392), .Y(n6715) );
  OAI21X1 U2327 ( .A(n5553), .B(n3388), .C(n6716), .Y(n9440) );
  NAND2X1 U2328 ( .A(arr[1138]), .B(n3392), .Y(n6716) );
  OAI21X1 U2329 ( .A(n5555), .B(n3388), .C(n6717), .Y(n9441) );
  NAND2X1 U2330 ( .A(arr[1139]), .B(n3392), .Y(n6717) );
  OAI21X1 U2331 ( .A(n5557), .B(n3388), .C(n6718), .Y(n9442) );
  NAND2X1 U2332 ( .A(arr[1140]), .B(n3392), .Y(n6718) );
  OAI21X1 U2333 ( .A(n5559), .B(n3387), .C(n6719), .Y(n9443) );
  NAND2X1 U2334 ( .A(arr[1141]), .B(n3392), .Y(n6719) );
  OAI21X1 U2335 ( .A(n5561), .B(n3387), .C(n6720), .Y(n9444) );
  NAND2X1 U2336 ( .A(arr[1142]), .B(n3392), .Y(n6720) );
  OAI21X1 U2337 ( .A(n5563), .B(n3387), .C(n6721), .Y(n9445) );
  NAND2X1 U2338 ( .A(arr[1143]), .B(n3392), .Y(n6721) );
  OAI21X1 U2339 ( .A(n5565), .B(n3387), .C(n6722), .Y(n9446) );
  NAND2X1 U2340 ( .A(arr[1144]), .B(n3392), .Y(n6722) );
  OAI21X1 U2341 ( .A(n5567), .B(n3387), .C(n6723), .Y(n9447) );
  NAND2X1 U2342 ( .A(arr[1145]), .B(n3392), .Y(n6723) );
  OAI21X1 U2343 ( .A(n5569), .B(n3387), .C(n6724), .Y(n9448) );
  NAND2X1 U2344 ( .A(arr[1146]), .B(n3390), .Y(n6724) );
  OAI21X1 U2345 ( .A(n5571), .B(n3387), .C(n6725), .Y(n9449) );
  NAND2X1 U2346 ( .A(arr[1147]), .B(n3390), .Y(n6725) );
  NAND2X1 U2347 ( .A(n6599), .B(n5703), .Y(n6684) );
  OAI21X1 U2349 ( .A(n5491), .B(n3381), .C(n6727), .Y(n9450) );
  NAND2X1 U2350 ( .A(arr[1148]), .B(n3384), .Y(n6727) );
  OAI21X1 U2351 ( .A(n5493), .B(n3381), .C(n6728), .Y(n9451) );
  NAND2X1 U2352 ( .A(arr[1149]), .B(n3384), .Y(n6728) );
  OAI21X1 U2353 ( .A(n5495), .B(n3381), .C(n6729), .Y(n9452) );
  NAND2X1 U2354 ( .A(arr[1150]), .B(n3384), .Y(n6729) );
  OAI21X1 U2355 ( .A(n5497), .B(n3381), .C(n6730), .Y(n9453) );
  NAND2X1 U2356 ( .A(arr[1151]), .B(n3384), .Y(n6730) );
  OAI21X1 U2357 ( .A(n5499), .B(n3381), .C(n6731), .Y(n9454) );
  NAND2X1 U2358 ( .A(arr[1152]), .B(n3384), .Y(n6731) );
  OAI21X1 U2359 ( .A(n5501), .B(n3382), .C(n6732), .Y(n9455) );
  NAND2X1 U2360 ( .A(arr[1153]), .B(n3384), .Y(n6732) );
  OAI21X1 U2361 ( .A(n5503), .B(n3382), .C(n6733), .Y(n9456) );
  NAND2X1 U2362 ( .A(arr[1154]), .B(n3384), .Y(n6733) );
  OAI21X1 U2363 ( .A(n5505), .B(n3382), .C(n6734), .Y(n9457) );
  NAND2X1 U2364 ( .A(arr[1155]), .B(n3384), .Y(n6734) );
  OAI21X1 U2365 ( .A(n5507), .B(n3381), .C(n6735), .Y(n9458) );
  NAND2X1 U2366 ( .A(arr[1156]), .B(n3384), .Y(n6735) );
  OAI21X1 U2367 ( .A(n5509), .B(n3382), .C(n6736), .Y(n9459) );
  NAND2X1 U2368 ( .A(arr[1157]), .B(n3384), .Y(n6736) );
  OAI21X1 U2369 ( .A(n5511), .B(n3383), .C(n6737), .Y(n9460) );
  NAND2X1 U2370 ( .A(arr[1158]), .B(n3384), .Y(n6737) );
  OAI21X1 U2371 ( .A(n5513), .B(n3383), .C(n6738), .Y(n9461) );
  NAND2X1 U2372 ( .A(arr[1159]), .B(n3384), .Y(n6738) );
  OAI21X1 U2373 ( .A(n5515), .B(n3383), .C(n6739), .Y(n9462) );
  NAND2X1 U2374 ( .A(arr[1160]), .B(n3384), .Y(n6739) );
  OAI21X1 U2375 ( .A(n5517), .B(n3382), .C(n6740), .Y(n9463) );
  NAND2X1 U2376 ( .A(arr[1161]), .B(n3385), .Y(n6740) );
  OAI21X1 U2377 ( .A(n5519), .B(n3384), .C(n6741), .Y(n9464) );
  NAND2X1 U2378 ( .A(arr[1162]), .B(n3385), .Y(n6741) );
  OAI21X1 U2379 ( .A(n5521), .B(n3384), .C(n6742), .Y(n9465) );
  NAND2X1 U2380 ( .A(arr[1163]), .B(n3385), .Y(n6742) );
  OAI21X1 U2381 ( .A(n5523), .B(n3383), .C(n6743), .Y(n9466) );
  NAND2X1 U2382 ( .A(arr[1164]), .B(n3385), .Y(n6743) );
  OAI21X1 U2383 ( .A(n5525), .B(n3383), .C(n6744), .Y(n9467) );
  NAND2X1 U2384 ( .A(arr[1165]), .B(n3385), .Y(n6744) );
  OAI21X1 U2385 ( .A(n5527), .B(n3383), .C(n6745), .Y(n9468) );
  NAND2X1 U2386 ( .A(arr[1166]), .B(n3385), .Y(n6745) );
  OAI21X1 U2387 ( .A(n5529), .B(n3383), .C(n6746), .Y(n9469) );
  NAND2X1 U2388 ( .A(arr[1167]), .B(n3385), .Y(n6746) );
  OAI21X1 U2389 ( .A(n5531), .B(n3383), .C(n6747), .Y(n9470) );
  NAND2X1 U2390 ( .A(arr[1168]), .B(n3385), .Y(n6747) );
  OAI21X1 U2391 ( .A(n5533), .B(n3383), .C(n6748), .Y(n9471) );
  NAND2X1 U2392 ( .A(arr[1169]), .B(n3385), .Y(n6748) );
  OAI21X1 U2393 ( .A(n5535), .B(n3383), .C(n6749), .Y(n9472) );
  NAND2X1 U2394 ( .A(arr[1170]), .B(n3385), .Y(n6749) );
  OAI21X1 U2395 ( .A(n5537), .B(n3383), .C(n6750), .Y(n9473) );
  NAND2X1 U2396 ( .A(arr[1171]), .B(n3385), .Y(n6750) );
  OAI21X1 U2397 ( .A(n5539), .B(n3383), .C(n6751), .Y(n9474) );
  NAND2X1 U2398 ( .A(arr[1172]), .B(n3385), .Y(n6751) );
  OAI21X1 U2399 ( .A(n5541), .B(n3383), .C(n6752), .Y(n9475) );
  NAND2X1 U2400 ( .A(arr[1173]), .B(n3385), .Y(n6752) );
  OAI21X1 U2401 ( .A(n5543), .B(n3382), .C(n6753), .Y(n9476) );
  NAND2X1 U2402 ( .A(arr[1174]), .B(n3385), .Y(n6753) );
  OAI21X1 U2403 ( .A(n5545), .B(n3382), .C(n6754), .Y(n9477) );
  NAND2X1 U2404 ( .A(arr[1175]), .B(n3385), .Y(n6754) );
  OAI21X1 U2405 ( .A(n5547), .B(n3382), .C(n6755), .Y(n9478) );
  NAND2X1 U2406 ( .A(arr[1176]), .B(n3385), .Y(n6755) );
  OAI21X1 U2407 ( .A(n5549), .B(n3382), .C(n6756), .Y(n9479) );
  NAND2X1 U2408 ( .A(arr[1177]), .B(n3385), .Y(n6756) );
  OAI21X1 U2409 ( .A(n5551), .B(n3382), .C(n6757), .Y(n9480) );
  NAND2X1 U2410 ( .A(arr[1178]), .B(n3386), .Y(n6757) );
  OAI21X1 U2411 ( .A(n5553), .B(n3382), .C(n6758), .Y(n9481) );
  NAND2X1 U2412 ( .A(arr[1179]), .B(n3386), .Y(n6758) );
  OAI21X1 U2413 ( .A(n5555), .B(n3382), .C(n6759), .Y(n9482) );
  NAND2X1 U2414 ( .A(arr[1180]), .B(n3386), .Y(n6759) );
  OAI21X1 U2415 ( .A(n5557), .B(n3382), .C(n6760), .Y(n9483) );
  NAND2X1 U2416 ( .A(arr[1181]), .B(n3386), .Y(n6760) );
  OAI21X1 U2417 ( .A(n5559), .B(n3381), .C(n6761), .Y(n9484) );
  NAND2X1 U2418 ( .A(arr[1182]), .B(n3386), .Y(n6761) );
  OAI21X1 U2419 ( .A(n5561), .B(n3381), .C(n6762), .Y(n9485) );
  NAND2X1 U2420 ( .A(arr[1183]), .B(n3386), .Y(n6762) );
  OAI21X1 U2421 ( .A(n5563), .B(n3381), .C(n6763), .Y(n9486) );
  NAND2X1 U2422 ( .A(arr[1184]), .B(n3386), .Y(n6763) );
  OAI21X1 U2423 ( .A(n5565), .B(n3381), .C(n6764), .Y(n9487) );
  NAND2X1 U2424 ( .A(arr[1185]), .B(n3386), .Y(n6764) );
  OAI21X1 U2425 ( .A(n5567), .B(n3381), .C(n6765), .Y(n9488) );
  NAND2X1 U2426 ( .A(arr[1186]), .B(n3386), .Y(n6765) );
  OAI21X1 U2427 ( .A(n5569), .B(n3381), .C(n6766), .Y(n9489) );
  NAND2X1 U2428 ( .A(arr[1187]), .B(n3384), .Y(n6766) );
  OAI21X1 U2429 ( .A(n5571), .B(n3381), .C(n6767), .Y(n9490) );
  NAND2X1 U2430 ( .A(arr[1188]), .B(n3384), .Y(n6767) );
  NAND2X1 U2431 ( .A(n6768), .B(n5573), .Y(n6726) );
  OAI21X1 U2432 ( .A(n5491), .B(n3375), .C(n6770), .Y(n9491) );
  NAND2X1 U2433 ( .A(arr[1189]), .B(n3378), .Y(n6770) );
  OAI21X1 U2434 ( .A(n5493), .B(n3375), .C(n6771), .Y(n9492) );
  NAND2X1 U2435 ( .A(arr[1190]), .B(n3378), .Y(n6771) );
  OAI21X1 U2436 ( .A(n5495), .B(n3375), .C(n6772), .Y(n9493) );
  NAND2X1 U2437 ( .A(arr[1191]), .B(n3378), .Y(n6772) );
  OAI21X1 U2438 ( .A(n5497), .B(n3375), .C(n6773), .Y(n9494) );
  NAND2X1 U2439 ( .A(arr[1192]), .B(n3378), .Y(n6773) );
  OAI21X1 U2440 ( .A(n5499), .B(n3375), .C(n6774), .Y(n9495) );
  NAND2X1 U2441 ( .A(arr[1193]), .B(n3378), .Y(n6774) );
  OAI21X1 U2442 ( .A(n5501), .B(n3376), .C(n6775), .Y(n9496) );
  NAND2X1 U2443 ( .A(arr[1194]), .B(n3378), .Y(n6775) );
  OAI21X1 U2444 ( .A(n5503), .B(n3376), .C(n6776), .Y(n9497) );
  NAND2X1 U2445 ( .A(arr[1195]), .B(n3378), .Y(n6776) );
  OAI21X1 U2446 ( .A(n5505), .B(n3376), .C(n6777), .Y(n9498) );
  NAND2X1 U2447 ( .A(arr[1196]), .B(n3378), .Y(n6777) );
  OAI21X1 U2448 ( .A(n5507), .B(n3375), .C(n6778), .Y(n9499) );
  NAND2X1 U2449 ( .A(arr[1197]), .B(n3378), .Y(n6778) );
  OAI21X1 U2450 ( .A(n5509), .B(n3376), .C(n6779), .Y(n9500) );
  NAND2X1 U2451 ( .A(arr[1198]), .B(n3378), .Y(n6779) );
  OAI21X1 U2452 ( .A(n5511), .B(n3377), .C(n6780), .Y(n9501) );
  NAND2X1 U2453 ( .A(arr[1199]), .B(n3378), .Y(n6780) );
  OAI21X1 U2454 ( .A(n5513), .B(n3377), .C(n6781), .Y(n9502) );
  NAND2X1 U2455 ( .A(arr[1200]), .B(n3378), .Y(n6781) );
  OAI21X1 U2456 ( .A(n5515), .B(n3377), .C(n6782), .Y(n9503) );
  NAND2X1 U2457 ( .A(arr[1201]), .B(n3378), .Y(n6782) );
  OAI21X1 U2458 ( .A(n5517), .B(n3376), .C(n6783), .Y(n9504) );
  NAND2X1 U2459 ( .A(arr[1202]), .B(n3379), .Y(n6783) );
  OAI21X1 U2460 ( .A(n5519), .B(n3378), .C(n6784), .Y(n9505) );
  NAND2X1 U2461 ( .A(arr[1203]), .B(n3379), .Y(n6784) );
  OAI21X1 U2462 ( .A(n5521), .B(n3378), .C(n6785), .Y(n9506) );
  NAND2X1 U2463 ( .A(arr[1204]), .B(n3379), .Y(n6785) );
  OAI21X1 U2464 ( .A(n5523), .B(n3377), .C(n6786), .Y(n9507) );
  NAND2X1 U2465 ( .A(arr[1205]), .B(n3379), .Y(n6786) );
  OAI21X1 U2466 ( .A(n5525), .B(n3377), .C(n6787), .Y(n9508) );
  NAND2X1 U2467 ( .A(arr[1206]), .B(n3379), .Y(n6787) );
  OAI21X1 U2468 ( .A(n5527), .B(n3377), .C(n6788), .Y(n9509) );
  NAND2X1 U2469 ( .A(arr[1207]), .B(n3379), .Y(n6788) );
  OAI21X1 U2470 ( .A(n5529), .B(n3377), .C(n6789), .Y(n9510) );
  NAND2X1 U2471 ( .A(arr[1208]), .B(n3379), .Y(n6789) );
  OAI21X1 U2472 ( .A(n5531), .B(n3377), .C(n6790), .Y(n9511) );
  NAND2X1 U2473 ( .A(arr[1209]), .B(n3379), .Y(n6790) );
  OAI21X1 U2474 ( .A(n5533), .B(n3377), .C(n6791), .Y(n9512) );
  NAND2X1 U2475 ( .A(arr[1210]), .B(n3379), .Y(n6791) );
  OAI21X1 U2476 ( .A(n5535), .B(n3377), .C(n6792), .Y(n9513) );
  NAND2X1 U2477 ( .A(arr[1211]), .B(n3379), .Y(n6792) );
  OAI21X1 U2478 ( .A(n5537), .B(n3377), .C(n6793), .Y(n9514) );
  NAND2X1 U2479 ( .A(arr[1212]), .B(n3379), .Y(n6793) );
  OAI21X1 U2480 ( .A(n5539), .B(n3377), .C(n6794), .Y(n9515) );
  NAND2X1 U2481 ( .A(arr[1213]), .B(n3379), .Y(n6794) );
  OAI21X1 U2482 ( .A(n5541), .B(n3377), .C(n6795), .Y(n9516) );
  NAND2X1 U2483 ( .A(arr[1214]), .B(n3379), .Y(n6795) );
  OAI21X1 U2484 ( .A(n5543), .B(n3376), .C(n6796), .Y(n9517) );
  NAND2X1 U2485 ( .A(arr[1215]), .B(n3379), .Y(n6796) );
  OAI21X1 U2486 ( .A(n5545), .B(n3376), .C(n6797), .Y(n9518) );
  NAND2X1 U2487 ( .A(arr[1216]), .B(n3379), .Y(n6797) );
  OAI21X1 U2488 ( .A(n5547), .B(n3376), .C(n6798), .Y(n9519) );
  NAND2X1 U2489 ( .A(arr[1217]), .B(n3379), .Y(n6798) );
  OAI21X1 U2490 ( .A(n5549), .B(n3376), .C(n6799), .Y(n9520) );
  NAND2X1 U2491 ( .A(arr[1218]), .B(n3379), .Y(n6799) );
  OAI21X1 U2492 ( .A(n5551), .B(n3376), .C(n6800), .Y(n9521) );
  NAND2X1 U2493 ( .A(arr[1219]), .B(n3380), .Y(n6800) );
  OAI21X1 U2494 ( .A(n5553), .B(n3376), .C(n6801), .Y(n9522) );
  NAND2X1 U2495 ( .A(arr[1220]), .B(n3380), .Y(n6801) );
  OAI21X1 U2496 ( .A(n5555), .B(n3376), .C(n6802), .Y(n9523) );
  NAND2X1 U2497 ( .A(arr[1221]), .B(n3380), .Y(n6802) );
  OAI21X1 U2498 ( .A(n5557), .B(n3376), .C(n6803), .Y(n9524) );
  NAND2X1 U2499 ( .A(arr[1222]), .B(n3380), .Y(n6803) );
  OAI21X1 U2500 ( .A(n5559), .B(n3375), .C(n6804), .Y(n9525) );
  NAND2X1 U2501 ( .A(arr[1223]), .B(n3380), .Y(n6804) );
  OAI21X1 U2502 ( .A(n5561), .B(n3375), .C(n6805), .Y(n9526) );
  NAND2X1 U2503 ( .A(arr[1224]), .B(n3380), .Y(n6805) );
  OAI21X1 U2504 ( .A(n5563), .B(n3375), .C(n6806), .Y(n9527) );
  NAND2X1 U2505 ( .A(arr[1225]), .B(n3380), .Y(n6806) );
  OAI21X1 U2506 ( .A(n5565), .B(n3375), .C(n6807), .Y(n9528) );
  NAND2X1 U2507 ( .A(arr[1226]), .B(n3380), .Y(n6807) );
  OAI21X1 U2508 ( .A(n5567), .B(n3375), .C(n6808), .Y(n9529) );
  NAND2X1 U2509 ( .A(arr[1227]), .B(n3380), .Y(n6808) );
  OAI21X1 U2510 ( .A(n5569), .B(n3375), .C(n6809), .Y(n9530) );
  NAND2X1 U2511 ( .A(arr[1228]), .B(n3378), .Y(n6809) );
  OAI21X1 U2512 ( .A(n5571), .B(n3375), .C(n6810), .Y(n9531) );
  NAND2X1 U2513 ( .A(arr[1229]), .B(n3378), .Y(n6810) );
  NAND2X1 U2514 ( .A(n6768), .B(n5617), .Y(n6769) );
  OAI21X1 U2515 ( .A(n5491), .B(n3369), .C(n6812), .Y(n9532) );
  NAND2X1 U2516 ( .A(arr[1230]), .B(n3372), .Y(n6812) );
  OAI21X1 U2517 ( .A(n5493), .B(n3369), .C(n6813), .Y(n9533) );
  NAND2X1 U2518 ( .A(arr[1231]), .B(n3372), .Y(n6813) );
  OAI21X1 U2519 ( .A(n5495), .B(n3369), .C(n6814), .Y(n9534) );
  NAND2X1 U2520 ( .A(arr[1232]), .B(n3372), .Y(n6814) );
  OAI21X1 U2521 ( .A(n5497), .B(n3369), .C(n6815), .Y(n9535) );
  NAND2X1 U2522 ( .A(arr[1233]), .B(n3372), .Y(n6815) );
  OAI21X1 U2523 ( .A(n5499), .B(n3369), .C(n6816), .Y(n9536) );
  NAND2X1 U2524 ( .A(arr[1234]), .B(n3372), .Y(n6816) );
  OAI21X1 U2525 ( .A(n5501), .B(n3370), .C(n6817), .Y(n9537) );
  NAND2X1 U2526 ( .A(arr[1235]), .B(n3372), .Y(n6817) );
  OAI21X1 U2527 ( .A(n5503), .B(n3370), .C(n6818), .Y(n9538) );
  NAND2X1 U2528 ( .A(arr[1236]), .B(n3372), .Y(n6818) );
  OAI21X1 U2529 ( .A(n5505), .B(n3370), .C(n6819), .Y(n9539) );
  NAND2X1 U2530 ( .A(arr[1237]), .B(n3372), .Y(n6819) );
  OAI21X1 U2531 ( .A(n5507), .B(n3369), .C(n6820), .Y(n9540) );
  NAND2X1 U2532 ( .A(arr[1238]), .B(n3372), .Y(n6820) );
  OAI21X1 U2533 ( .A(n5509), .B(n3370), .C(n6821), .Y(n9541) );
  NAND2X1 U2534 ( .A(arr[1239]), .B(n3372), .Y(n6821) );
  OAI21X1 U2535 ( .A(n5511), .B(n3371), .C(n6822), .Y(n9542) );
  NAND2X1 U2536 ( .A(arr[1240]), .B(n3372), .Y(n6822) );
  OAI21X1 U2537 ( .A(n5513), .B(n3371), .C(n6823), .Y(n9543) );
  NAND2X1 U2538 ( .A(arr[1241]), .B(n3372), .Y(n6823) );
  OAI21X1 U2539 ( .A(n5515), .B(n3371), .C(n6824), .Y(n9544) );
  NAND2X1 U2540 ( .A(arr[1242]), .B(n3372), .Y(n6824) );
  OAI21X1 U2541 ( .A(n5517), .B(n3370), .C(n6825), .Y(n9545) );
  NAND2X1 U2542 ( .A(arr[1243]), .B(n3373), .Y(n6825) );
  OAI21X1 U2543 ( .A(n5519), .B(n3372), .C(n6826), .Y(n9546) );
  NAND2X1 U2544 ( .A(arr[1244]), .B(n3373), .Y(n6826) );
  OAI21X1 U2545 ( .A(n5521), .B(n3372), .C(n6827), .Y(n9547) );
  NAND2X1 U2546 ( .A(arr[1245]), .B(n3373), .Y(n6827) );
  OAI21X1 U2547 ( .A(n5523), .B(n3371), .C(n6828), .Y(n9548) );
  NAND2X1 U2548 ( .A(arr[1246]), .B(n3373), .Y(n6828) );
  OAI21X1 U2549 ( .A(n5525), .B(n3371), .C(n6829), .Y(n9549) );
  NAND2X1 U2550 ( .A(arr[1247]), .B(n3373), .Y(n6829) );
  OAI21X1 U2551 ( .A(n5527), .B(n3371), .C(n6830), .Y(n9550) );
  NAND2X1 U2552 ( .A(arr[1248]), .B(n3373), .Y(n6830) );
  OAI21X1 U2553 ( .A(n5529), .B(n3371), .C(n6831), .Y(n9551) );
  NAND2X1 U2554 ( .A(arr[1249]), .B(n3373), .Y(n6831) );
  OAI21X1 U2555 ( .A(n5531), .B(n3371), .C(n6832), .Y(n9552) );
  NAND2X1 U2556 ( .A(arr[1250]), .B(n3373), .Y(n6832) );
  OAI21X1 U2557 ( .A(n5533), .B(n3371), .C(n6833), .Y(n9553) );
  NAND2X1 U2558 ( .A(arr[1251]), .B(n3373), .Y(n6833) );
  OAI21X1 U2559 ( .A(n5535), .B(n3371), .C(n6834), .Y(n9554) );
  NAND2X1 U2560 ( .A(arr[1252]), .B(n3373), .Y(n6834) );
  OAI21X1 U2561 ( .A(n5537), .B(n3371), .C(n6835), .Y(n9555) );
  NAND2X1 U2562 ( .A(arr[1253]), .B(n3373), .Y(n6835) );
  OAI21X1 U2563 ( .A(n5539), .B(n3371), .C(n6836), .Y(n9556) );
  NAND2X1 U2564 ( .A(arr[1254]), .B(n3373), .Y(n6836) );
  OAI21X1 U2565 ( .A(n5541), .B(n3371), .C(n6837), .Y(n9557) );
  NAND2X1 U2566 ( .A(arr[1255]), .B(n3373), .Y(n6837) );
  OAI21X1 U2567 ( .A(n5543), .B(n3370), .C(n6838), .Y(n9558) );
  NAND2X1 U2568 ( .A(arr[1256]), .B(n3373), .Y(n6838) );
  OAI21X1 U2569 ( .A(n5545), .B(n3370), .C(n6839), .Y(n9559) );
  NAND2X1 U2570 ( .A(arr[1257]), .B(n3373), .Y(n6839) );
  OAI21X1 U2571 ( .A(n5547), .B(n3370), .C(n6840), .Y(n9560) );
  NAND2X1 U2572 ( .A(arr[1258]), .B(n3373), .Y(n6840) );
  OAI21X1 U2573 ( .A(n5549), .B(n3370), .C(n6841), .Y(n9561) );
  NAND2X1 U2574 ( .A(arr[1259]), .B(n3373), .Y(n6841) );
  OAI21X1 U2575 ( .A(n5551), .B(n3370), .C(n6842), .Y(n9562) );
  NAND2X1 U2576 ( .A(arr[1260]), .B(n3374), .Y(n6842) );
  OAI21X1 U2577 ( .A(n5553), .B(n3370), .C(n6843), .Y(n9563) );
  NAND2X1 U2578 ( .A(arr[1261]), .B(n3374), .Y(n6843) );
  OAI21X1 U2579 ( .A(n5555), .B(n3370), .C(n6844), .Y(n9564) );
  NAND2X1 U2580 ( .A(arr[1262]), .B(n3374), .Y(n6844) );
  OAI21X1 U2581 ( .A(n5557), .B(n3370), .C(n6845), .Y(n9565) );
  NAND2X1 U2582 ( .A(arr[1263]), .B(n3374), .Y(n6845) );
  OAI21X1 U2583 ( .A(n5559), .B(n3369), .C(n6846), .Y(n9566) );
  NAND2X1 U2584 ( .A(arr[1264]), .B(n3374), .Y(n6846) );
  OAI21X1 U2585 ( .A(n5561), .B(n3369), .C(n6847), .Y(n9567) );
  NAND2X1 U2586 ( .A(arr[1265]), .B(n3374), .Y(n6847) );
  OAI21X1 U2587 ( .A(n5563), .B(n3369), .C(n6848), .Y(n9568) );
  NAND2X1 U2588 ( .A(arr[1266]), .B(n3374), .Y(n6848) );
  OAI21X1 U2589 ( .A(n5565), .B(n3369), .C(n6849), .Y(n9569) );
  NAND2X1 U2590 ( .A(arr[1267]), .B(n3374), .Y(n6849) );
  OAI21X1 U2591 ( .A(n5567), .B(n3369), .C(n6850), .Y(n9570) );
  NAND2X1 U2592 ( .A(arr[1268]), .B(n3374), .Y(n6850) );
  OAI21X1 U2593 ( .A(n5569), .B(n3369), .C(n6851), .Y(n9571) );
  NAND2X1 U2594 ( .A(arr[1269]), .B(n3372), .Y(n6851) );
  OAI21X1 U2595 ( .A(n5571), .B(n3369), .C(n6852), .Y(n9572) );
  NAND2X1 U2596 ( .A(arr[1270]), .B(n3372), .Y(n6852) );
  NAND2X1 U2597 ( .A(n6768), .B(n5660), .Y(n6811) );
  OAI21X1 U2598 ( .A(n5491), .B(n3363), .C(n6854), .Y(n9573) );
  NAND2X1 U2599 ( .A(arr[1271]), .B(n3366), .Y(n6854) );
  OAI21X1 U2600 ( .A(n5493), .B(n3363), .C(n6855), .Y(n9574) );
  NAND2X1 U2601 ( .A(arr[1272]), .B(n3366), .Y(n6855) );
  OAI21X1 U2602 ( .A(n5495), .B(n3363), .C(n6856), .Y(n9575) );
  NAND2X1 U2603 ( .A(arr[1273]), .B(n3366), .Y(n6856) );
  OAI21X1 U2604 ( .A(n5497), .B(n3363), .C(n6857), .Y(n9576) );
  NAND2X1 U2605 ( .A(arr[1274]), .B(n3366), .Y(n6857) );
  OAI21X1 U2606 ( .A(n5499), .B(n3363), .C(n6858), .Y(n9577) );
  NAND2X1 U2607 ( .A(arr[1275]), .B(n3366), .Y(n6858) );
  OAI21X1 U2608 ( .A(n5501), .B(n3364), .C(n6859), .Y(n9578) );
  NAND2X1 U2609 ( .A(arr[1276]), .B(n3366), .Y(n6859) );
  OAI21X1 U2610 ( .A(n5503), .B(n3364), .C(n6860), .Y(n9579) );
  NAND2X1 U2611 ( .A(arr[1277]), .B(n3366), .Y(n6860) );
  OAI21X1 U2612 ( .A(n5505), .B(n3364), .C(n6861), .Y(n9580) );
  NAND2X1 U2613 ( .A(arr[1278]), .B(n3366), .Y(n6861) );
  OAI21X1 U2614 ( .A(n5507), .B(n3363), .C(n6862), .Y(n9581) );
  NAND2X1 U2615 ( .A(arr[1279]), .B(n3366), .Y(n6862) );
  OAI21X1 U2616 ( .A(n5509), .B(n3364), .C(n6863), .Y(n9582) );
  NAND2X1 U2617 ( .A(arr[1280]), .B(n3366), .Y(n6863) );
  OAI21X1 U2618 ( .A(n5511), .B(n3365), .C(n6864), .Y(n9583) );
  NAND2X1 U2619 ( .A(arr[1281]), .B(n3366), .Y(n6864) );
  OAI21X1 U2620 ( .A(n5513), .B(n3365), .C(n6865), .Y(n9584) );
  NAND2X1 U2621 ( .A(arr[1282]), .B(n3366), .Y(n6865) );
  OAI21X1 U2622 ( .A(n5515), .B(n3365), .C(n6866), .Y(n9585) );
  NAND2X1 U2623 ( .A(arr[1283]), .B(n3366), .Y(n6866) );
  OAI21X1 U2624 ( .A(n5517), .B(n3364), .C(n6867), .Y(n9586) );
  NAND2X1 U2625 ( .A(arr[1284]), .B(n3367), .Y(n6867) );
  OAI21X1 U2626 ( .A(n5519), .B(n3366), .C(n6868), .Y(n9587) );
  NAND2X1 U2627 ( .A(arr[1285]), .B(n3367), .Y(n6868) );
  OAI21X1 U2628 ( .A(n5521), .B(n3366), .C(n6869), .Y(n9588) );
  NAND2X1 U2629 ( .A(arr[1286]), .B(n3367), .Y(n6869) );
  OAI21X1 U2630 ( .A(n5523), .B(n3365), .C(n6870), .Y(n9589) );
  NAND2X1 U2631 ( .A(arr[1287]), .B(n3367), .Y(n6870) );
  OAI21X1 U2632 ( .A(n5525), .B(n3365), .C(n6871), .Y(n9590) );
  NAND2X1 U2633 ( .A(arr[1288]), .B(n3367), .Y(n6871) );
  OAI21X1 U2634 ( .A(n5527), .B(n3365), .C(n6872), .Y(n9591) );
  NAND2X1 U2635 ( .A(arr[1289]), .B(n3367), .Y(n6872) );
  OAI21X1 U2636 ( .A(n5529), .B(n3365), .C(n6873), .Y(n9592) );
  NAND2X1 U2637 ( .A(arr[1290]), .B(n3367), .Y(n6873) );
  OAI21X1 U2638 ( .A(n5531), .B(n3365), .C(n6874), .Y(n9593) );
  NAND2X1 U2639 ( .A(arr[1291]), .B(n3367), .Y(n6874) );
  OAI21X1 U2640 ( .A(n5533), .B(n3365), .C(n6875), .Y(n9594) );
  NAND2X1 U2641 ( .A(arr[1292]), .B(n3367), .Y(n6875) );
  OAI21X1 U2642 ( .A(n5535), .B(n3365), .C(n6876), .Y(n9595) );
  NAND2X1 U2643 ( .A(arr[1293]), .B(n3367), .Y(n6876) );
  OAI21X1 U2644 ( .A(n5537), .B(n3365), .C(n6877), .Y(n9596) );
  NAND2X1 U2645 ( .A(arr[1294]), .B(n3367), .Y(n6877) );
  OAI21X1 U2646 ( .A(n5539), .B(n3365), .C(n6878), .Y(n9597) );
  NAND2X1 U2647 ( .A(arr[1295]), .B(n3367), .Y(n6878) );
  OAI21X1 U2648 ( .A(n5541), .B(n3365), .C(n6879), .Y(n9598) );
  NAND2X1 U2649 ( .A(arr[1296]), .B(n3367), .Y(n6879) );
  OAI21X1 U2650 ( .A(n5543), .B(n3364), .C(n6880), .Y(n9599) );
  NAND2X1 U2651 ( .A(arr[1297]), .B(n3367), .Y(n6880) );
  OAI21X1 U2652 ( .A(n5545), .B(n3364), .C(n6881), .Y(n9600) );
  NAND2X1 U2653 ( .A(arr[1298]), .B(n3367), .Y(n6881) );
  OAI21X1 U2654 ( .A(n5547), .B(n3364), .C(n6882), .Y(n9601) );
  NAND2X1 U2655 ( .A(arr[1299]), .B(n3367), .Y(n6882) );
  OAI21X1 U2656 ( .A(n5549), .B(n3364), .C(n6883), .Y(n9602) );
  NAND2X1 U2657 ( .A(arr[1300]), .B(n3367), .Y(n6883) );
  OAI21X1 U2658 ( .A(n5551), .B(n3364), .C(n6884), .Y(n9603) );
  NAND2X1 U2659 ( .A(arr[1301]), .B(n3368), .Y(n6884) );
  OAI21X1 U2660 ( .A(n5553), .B(n3364), .C(n6885), .Y(n9604) );
  NAND2X1 U2661 ( .A(arr[1302]), .B(n3368), .Y(n6885) );
  OAI21X1 U2662 ( .A(n5555), .B(n3364), .C(n6886), .Y(n9605) );
  NAND2X1 U2663 ( .A(arr[1303]), .B(n3368), .Y(n6886) );
  OAI21X1 U2664 ( .A(n5557), .B(n3364), .C(n6887), .Y(n9606) );
  NAND2X1 U2665 ( .A(arr[1304]), .B(n3368), .Y(n6887) );
  OAI21X1 U2666 ( .A(n5559), .B(n3363), .C(n6888), .Y(n9607) );
  NAND2X1 U2667 ( .A(arr[1305]), .B(n3368), .Y(n6888) );
  OAI21X1 U2668 ( .A(n5561), .B(n3363), .C(n6889), .Y(n9608) );
  NAND2X1 U2669 ( .A(arr[1306]), .B(n3368), .Y(n6889) );
  OAI21X1 U2670 ( .A(n5563), .B(n3363), .C(n6890), .Y(n9609) );
  NAND2X1 U2671 ( .A(arr[1307]), .B(n3368), .Y(n6890) );
  OAI21X1 U2672 ( .A(n5565), .B(n3363), .C(n6891), .Y(n9610) );
  NAND2X1 U2673 ( .A(arr[1308]), .B(n3368), .Y(n6891) );
  OAI21X1 U2674 ( .A(n5567), .B(n3363), .C(n6892), .Y(n9611) );
  NAND2X1 U2675 ( .A(arr[1309]), .B(n3368), .Y(n6892) );
  OAI21X1 U2676 ( .A(n5569), .B(n3363), .C(n6893), .Y(n9612) );
  NAND2X1 U2677 ( .A(arr[1310]), .B(n3366), .Y(n6893) );
  OAI21X1 U2678 ( .A(n5571), .B(n3363), .C(n6894), .Y(n9613) );
  NAND2X1 U2679 ( .A(arr[1311]), .B(n3366), .Y(n6894) );
  NAND2X1 U2680 ( .A(n6768), .B(n5703), .Y(n6853) );
  AND2X1 U2682 ( .A(wr_ptr[4]), .B(n6216), .Y(n6387) );
  AND2X1 U2683 ( .A(n6895), .B(n6896), .Y(n6216) );
  OAI21X1 U2684 ( .A(n5491), .B(n3357), .C(n6898), .Y(n9614) );
  NAND2X1 U2685 ( .A(arr[1312]), .B(n3360), .Y(n6898) );
  OAI21X1 U2686 ( .A(n5493), .B(n3357), .C(n6899), .Y(n9615) );
  NAND2X1 U2687 ( .A(arr[1313]), .B(n3360), .Y(n6899) );
  OAI21X1 U2688 ( .A(n5495), .B(n3357), .C(n6900), .Y(n9616) );
  NAND2X1 U2689 ( .A(arr[1314]), .B(n3360), .Y(n6900) );
  OAI21X1 U2690 ( .A(n5497), .B(n3357), .C(n6901), .Y(n9617) );
  NAND2X1 U2691 ( .A(arr[1315]), .B(n3360), .Y(n6901) );
  OAI21X1 U2692 ( .A(n5499), .B(n3357), .C(n6902), .Y(n9618) );
  NAND2X1 U2693 ( .A(arr[1316]), .B(n3360), .Y(n6902) );
  OAI21X1 U2694 ( .A(n5501), .B(n3358), .C(n6903), .Y(n9619) );
  NAND2X1 U2695 ( .A(arr[1317]), .B(n3360), .Y(n6903) );
  OAI21X1 U2696 ( .A(n5503), .B(n3358), .C(n6904), .Y(n9620) );
  NAND2X1 U2697 ( .A(arr[1318]), .B(n3360), .Y(n6904) );
  OAI21X1 U2698 ( .A(n5505), .B(n3358), .C(n6905), .Y(n9621) );
  NAND2X1 U2699 ( .A(arr[1319]), .B(n3360), .Y(n6905) );
  OAI21X1 U2700 ( .A(n5507), .B(n3357), .C(n6906), .Y(n9622) );
  NAND2X1 U2701 ( .A(arr[1320]), .B(n3360), .Y(n6906) );
  OAI21X1 U2702 ( .A(n5509), .B(n3358), .C(n6907), .Y(n9623) );
  NAND2X1 U2703 ( .A(arr[1321]), .B(n3360), .Y(n6907) );
  OAI21X1 U2704 ( .A(n5511), .B(n3359), .C(n6908), .Y(n9624) );
  NAND2X1 U2705 ( .A(arr[1322]), .B(n3360), .Y(n6908) );
  OAI21X1 U2706 ( .A(n5513), .B(n3359), .C(n6909), .Y(n9625) );
  NAND2X1 U2707 ( .A(arr[1323]), .B(n3360), .Y(n6909) );
  OAI21X1 U2708 ( .A(n5515), .B(n3359), .C(n6910), .Y(n9626) );
  NAND2X1 U2709 ( .A(arr[1324]), .B(n3360), .Y(n6910) );
  OAI21X1 U2710 ( .A(n5517), .B(n3358), .C(n6911), .Y(n9627) );
  NAND2X1 U2711 ( .A(arr[1325]), .B(n3361), .Y(n6911) );
  OAI21X1 U2712 ( .A(n5519), .B(n3360), .C(n6912), .Y(n9628) );
  NAND2X1 U2713 ( .A(arr[1326]), .B(n3361), .Y(n6912) );
  OAI21X1 U2714 ( .A(n5521), .B(n3360), .C(n6913), .Y(n9629) );
  NAND2X1 U2715 ( .A(arr[1327]), .B(n3361), .Y(n6913) );
  OAI21X1 U2716 ( .A(n5523), .B(n3359), .C(n6914), .Y(n9630) );
  NAND2X1 U2717 ( .A(arr[1328]), .B(n3361), .Y(n6914) );
  OAI21X1 U2718 ( .A(n5525), .B(n3359), .C(n6915), .Y(n9631) );
  NAND2X1 U2719 ( .A(arr[1329]), .B(n3361), .Y(n6915) );
  OAI21X1 U2720 ( .A(n5527), .B(n3359), .C(n6916), .Y(n9632) );
  NAND2X1 U2721 ( .A(arr[1330]), .B(n3361), .Y(n6916) );
  OAI21X1 U2722 ( .A(n5529), .B(n3359), .C(n6917), .Y(n9633) );
  NAND2X1 U2723 ( .A(arr[1331]), .B(n3361), .Y(n6917) );
  OAI21X1 U2724 ( .A(n5531), .B(n3359), .C(n6918), .Y(n9634) );
  NAND2X1 U2725 ( .A(arr[1332]), .B(n3361), .Y(n6918) );
  OAI21X1 U2726 ( .A(n5533), .B(n3359), .C(n6919), .Y(n9635) );
  NAND2X1 U2727 ( .A(arr[1333]), .B(n3361), .Y(n6919) );
  OAI21X1 U2728 ( .A(n5535), .B(n3359), .C(n6920), .Y(n9636) );
  NAND2X1 U2729 ( .A(arr[1334]), .B(n3361), .Y(n6920) );
  OAI21X1 U2730 ( .A(n5537), .B(n3359), .C(n6921), .Y(n9637) );
  NAND2X1 U2731 ( .A(arr[1335]), .B(n3361), .Y(n6921) );
  OAI21X1 U2732 ( .A(n5539), .B(n3359), .C(n6922), .Y(n9638) );
  NAND2X1 U2733 ( .A(arr[1336]), .B(n3361), .Y(n6922) );
  OAI21X1 U2734 ( .A(n5541), .B(n3359), .C(n6923), .Y(n9639) );
  NAND2X1 U2735 ( .A(arr[1337]), .B(n3361), .Y(n6923) );
  OAI21X1 U2736 ( .A(n5543), .B(n3358), .C(n6924), .Y(n9640) );
  NAND2X1 U2737 ( .A(arr[1338]), .B(n3361), .Y(n6924) );
  OAI21X1 U2738 ( .A(n5545), .B(n3358), .C(n6925), .Y(n9641) );
  NAND2X1 U2739 ( .A(arr[1339]), .B(n3361), .Y(n6925) );
  OAI21X1 U2740 ( .A(n5547), .B(n3358), .C(n6926), .Y(n9642) );
  NAND2X1 U2741 ( .A(arr[1340]), .B(n3361), .Y(n6926) );
  OAI21X1 U2742 ( .A(n5549), .B(n3358), .C(n6927), .Y(n9643) );
  NAND2X1 U2743 ( .A(arr[1341]), .B(n3361), .Y(n6927) );
  OAI21X1 U2744 ( .A(n5551), .B(n3358), .C(n6928), .Y(n9644) );
  NAND2X1 U2745 ( .A(arr[1342]), .B(n3362), .Y(n6928) );
  OAI21X1 U2746 ( .A(n5553), .B(n3358), .C(n6929), .Y(n9645) );
  NAND2X1 U2747 ( .A(arr[1343]), .B(n3362), .Y(n6929) );
  OAI21X1 U2748 ( .A(n5555), .B(n3358), .C(n6930), .Y(n9646) );
  NAND2X1 U2749 ( .A(arr[1344]), .B(n3362), .Y(n6930) );
  OAI21X1 U2750 ( .A(n5557), .B(n3358), .C(n6931), .Y(n9647) );
  NAND2X1 U2751 ( .A(arr[1345]), .B(n3362), .Y(n6931) );
  OAI21X1 U2752 ( .A(n5559), .B(n3357), .C(n6932), .Y(n9648) );
  NAND2X1 U2753 ( .A(arr[1346]), .B(n3362), .Y(n6932) );
  OAI21X1 U2754 ( .A(n5561), .B(n3357), .C(n6933), .Y(n9649) );
  NAND2X1 U2755 ( .A(arr[1347]), .B(n3362), .Y(n6933) );
  OAI21X1 U2756 ( .A(n5563), .B(n3357), .C(n6934), .Y(n9650) );
  NAND2X1 U2757 ( .A(arr[1348]), .B(n3362), .Y(n6934) );
  OAI21X1 U2758 ( .A(n5565), .B(n3357), .C(n6935), .Y(n9651) );
  NAND2X1 U2759 ( .A(arr[1349]), .B(n3362), .Y(n6935) );
  OAI21X1 U2760 ( .A(n5567), .B(n3357), .C(n6936), .Y(n9652) );
  NAND2X1 U2761 ( .A(arr[1350]), .B(n3362), .Y(n6936) );
  OAI21X1 U2762 ( .A(n5569), .B(n3357), .C(n6937), .Y(n9653) );
  NAND2X1 U2763 ( .A(arr[1351]), .B(n3360), .Y(n6937) );
  OAI21X1 U2764 ( .A(n5571), .B(n3357), .C(n6938), .Y(n9654) );
  NAND2X1 U2765 ( .A(arr[1352]), .B(n3360), .Y(n6938) );
  NAND2X1 U2766 ( .A(n6939), .B(n5573), .Y(n6897) );
  OAI21X1 U2767 ( .A(n5491), .B(n3351), .C(n6941), .Y(n9655) );
  NAND2X1 U2768 ( .A(arr[1353]), .B(n3354), .Y(n6941) );
  OAI21X1 U2769 ( .A(n5493), .B(n3351), .C(n6942), .Y(n9656) );
  NAND2X1 U2770 ( .A(arr[1354]), .B(n3354), .Y(n6942) );
  OAI21X1 U2771 ( .A(n5495), .B(n3351), .C(n6943), .Y(n9657) );
  NAND2X1 U2772 ( .A(arr[1355]), .B(n3354), .Y(n6943) );
  OAI21X1 U2773 ( .A(n5497), .B(n3351), .C(n6944), .Y(n9658) );
  NAND2X1 U2774 ( .A(arr[1356]), .B(n3354), .Y(n6944) );
  OAI21X1 U2775 ( .A(n5499), .B(n3351), .C(n6945), .Y(n9659) );
  NAND2X1 U2776 ( .A(arr[1357]), .B(n3354), .Y(n6945) );
  OAI21X1 U2777 ( .A(n5501), .B(n3352), .C(n6946), .Y(n9660) );
  NAND2X1 U2778 ( .A(arr[1358]), .B(n3354), .Y(n6946) );
  OAI21X1 U2779 ( .A(n5503), .B(n3352), .C(n6947), .Y(n9661) );
  NAND2X1 U2780 ( .A(arr[1359]), .B(n3354), .Y(n6947) );
  OAI21X1 U2781 ( .A(n5505), .B(n3352), .C(n6948), .Y(n9662) );
  NAND2X1 U2782 ( .A(arr[1360]), .B(n3354), .Y(n6948) );
  OAI21X1 U2783 ( .A(n5507), .B(n3351), .C(n6949), .Y(n9663) );
  NAND2X1 U2784 ( .A(arr[1361]), .B(n3354), .Y(n6949) );
  OAI21X1 U2785 ( .A(n5509), .B(n3352), .C(n6950), .Y(n9664) );
  NAND2X1 U2786 ( .A(arr[1362]), .B(n3354), .Y(n6950) );
  OAI21X1 U2787 ( .A(n5511), .B(n3353), .C(n6951), .Y(n9665) );
  NAND2X1 U2788 ( .A(arr[1363]), .B(n3354), .Y(n6951) );
  OAI21X1 U2789 ( .A(n5513), .B(n3353), .C(n6952), .Y(n9666) );
  NAND2X1 U2790 ( .A(arr[1364]), .B(n3354), .Y(n6952) );
  OAI21X1 U2791 ( .A(n5515), .B(n3353), .C(n6953), .Y(n9667) );
  NAND2X1 U2792 ( .A(arr[1365]), .B(n3354), .Y(n6953) );
  OAI21X1 U2793 ( .A(n5517), .B(n3352), .C(n6954), .Y(n9668) );
  NAND2X1 U2794 ( .A(arr[1366]), .B(n3355), .Y(n6954) );
  OAI21X1 U2795 ( .A(n5519), .B(n3354), .C(n6955), .Y(n9669) );
  NAND2X1 U2796 ( .A(arr[1367]), .B(n3355), .Y(n6955) );
  OAI21X1 U2797 ( .A(n5521), .B(n3354), .C(n6956), .Y(n9670) );
  NAND2X1 U2798 ( .A(arr[1368]), .B(n3355), .Y(n6956) );
  OAI21X1 U2799 ( .A(n5523), .B(n3353), .C(n6957), .Y(n9671) );
  NAND2X1 U2800 ( .A(arr[1369]), .B(n3355), .Y(n6957) );
  OAI21X1 U2801 ( .A(n5525), .B(n3353), .C(n6958), .Y(n9672) );
  NAND2X1 U2802 ( .A(arr[1370]), .B(n3355), .Y(n6958) );
  OAI21X1 U2803 ( .A(n5527), .B(n3353), .C(n6959), .Y(n9673) );
  NAND2X1 U2804 ( .A(arr[1371]), .B(n3355), .Y(n6959) );
  OAI21X1 U2805 ( .A(n5529), .B(n3353), .C(n6960), .Y(n9674) );
  NAND2X1 U2806 ( .A(arr[1372]), .B(n3355), .Y(n6960) );
  OAI21X1 U2807 ( .A(n5531), .B(n3353), .C(n6961), .Y(n9675) );
  NAND2X1 U2808 ( .A(arr[1373]), .B(n3355), .Y(n6961) );
  OAI21X1 U2809 ( .A(n5533), .B(n3353), .C(n6962), .Y(n9676) );
  NAND2X1 U2810 ( .A(arr[1374]), .B(n3355), .Y(n6962) );
  OAI21X1 U2811 ( .A(n5535), .B(n3353), .C(n6963), .Y(n9677) );
  NAND2X1 U2812 ( .A(arr[1375]), .B(n3355), .Y(n6963) );
  OAI21X1 U2813 ( .A(n5537), .B(n3353), .C(n6964), .Y(n9678) );
  NAND2X1 U2814 ( .A(arr[1376]), .B(n3355), .Y(n6964) );
  OAI21X1 U2815 ( .A(n5539), .B(n3353), .C(n6965), .Y(n9679) );
  NAND2X1 U2816 ( .A(arr[1377]), .B(n3355), .Y(n6965) );
  OAI21X1 U2817 ( .A(n5541), .B(n3353), .C(n6966), .Y(n9680) );
  NAND2X1 U2818 ( .A(arr[1378]), .B(n3355), .Y(n6966) );
  OAI21X1 U2819 ( .A(n5543), .B(n3352), .C(n6967), .Y(n9681) );
  NAND2X1 U2820 ( .A(arr[1379]), .B(n3355), .Y(n6967) );
  OAI21X1 U2821 ( .A(n5545), .B(n3352), .C(n6968), .Y(n9682) );
  NAND2X1 U2822 ( .A(arr[1380]), .B(n3355), .Y(n6968) );
  OAI21X1 U2823 ( .A(n5547), .B(n3352), .C(n6969), .Y(n9683) );
  NAND2X1 U2824 ( .A(arr[1381]), .B(n3355), .Y(n6969) );
  OAI21X1 U2825 ( .A(n5549), .B(n3352), .C(n6970), .Y(n9684) );
  NAND2X1 U2826 ( .A(arr[1382]), .B(n3355), .Y(n6970) );
  OAI21X1 U2827 ( .A(n5551), .B(n3352), .C(n6971), .Y(n9685) );
  NAND2X1 U2828 ( .A(arr[1383]), .B(n3356), .Y(n6971) );
  OAI21X1 U2829 ( .A(n5553), .B(n3352), .C(n6972), .Y(n9686) );
  NAND2X1 U2830 ( .A(arr[1384]), .B(n3356), .Y(n6972) );
  OAI21X1 U2831 ( .A(n5555), .B(n3352), .C(n6973), .Y(n9687) );
  NAND2X1 U2832 ( .A(arr[1385]), .B(n3356), .Y(n6973) );
  OAI21X1 U2833 ( .A(n5557), .B(n3352), .C(n6974), .Y(n9688) );
  NAND2X1 U2834 ( .A(arr[1386]), .B(n3356), .Y(n6974) );
  OAI21X1 U2835 ( .A(n5559), .B(n3351), .C(n6975), .Y(n9689) );
  NAND2X1 U2836 ( .A(arr[1387]), .B(n3356), .Y(n6975) );
  OAI21X1 U2837 ( .A(n5561), .B(n3351), .C(n6976), .Y(n9690) );
  NAND2X1 U2838 ( .A(arr[1388]), .B(n3356), .Y(n6976) );
  OAI21X1 U2839 ( .A(n5563), .B(n3351), .C(n6977), .Y(n9691) );
  NAND2X1 U2840 ( .A(arr[1389]), .B(n3356), .Y(n6977) );
  OAI21X1 U2841 ( .A(n5565), .B(n3351), .C(n6978), .Y(n9692) );
  NAND2X1 U2842 ( .A(arr[1390]), .B(n3356), .Y(n6978) );
  OAI21X1 U2843 ( .A(n5567), .B(n3351), .C(n6979), .Y(n9693) );
  NAND2X1 U2844 ( .A(arr[1391]), .B(n3356), .Y(n6979) );
  OAI21X1 U2845 ( .A(n5569), .B(n3351), .C(n6980), .Y(n9694) );
  NAND2X1 U2846 ( .A(arr[1392]), .B(n3354), .Y(n6980) );
  OAI21X1 U2847 ( .A(n5571), .B(n3356), .C(n6981), .Y(n9695) );
  NAND2X1 U2848 ( .A(arr[1393]), .B(n3354), .Y(n6981) );
  NAND2X1 U2849 ( .A(n6939), .B(n5617), .Y(n6940) );
  OAI21X1 U2850 ( .A(n5491), .B(n3345), .C(n6983), .Y(n9696) );
  NAND2X1 U2851 ( .A(arr[1394]), .B(n3348), .Y(n6983) );
  OAI21X1 U2852 ( .A(n5493), .B(n3345), .C(n6984), .Y(n9697) );
  NAND2X1 U2853 ( .A(arr[1395]), .B(n3348), .Y(n6984) );
  OAI21X1 U2854 ( .A(n5495), .B(n3345), .C(n6985), .Y(n9698) );
  NAND2X1 U2855 ( .A(arr[1396]), .B(n3348), .Y(n6985) );
  OAI21X1 U2856 ( .A(n5497), .B(n3345), .C(n6986), .Y(n9699) );
  NAND2X1 U2857 ( .A(arr[1397]), .B(n3348), .Y(n6986) );
  OAI21X1 U2858 ( .A(n5499), .B(n3345), .C(n6987), .Y(n9700) );
  NAND2X1 U2859 ( .A(arr[1398]), .B(n3348), .Y(n6987) );
  OAI21X1 U2860 ( .A(n5501), .B(n3346), .C(n6988), .Y(n9701) );
  NAND2X1 U2861 ( .A(arr[1399]), .B(n3348), .Y(n6988) );
  OAI21X1 U2862 ( .A(n5503), .B(n3346), .C(n6989), .Y(n9702) );
  NAND2X1 U2863 ( .A(arr[1400]), .B(n3348), .Y(n6989) );
  OAI21X1 U2864 ( .A(n5505), .B(n3346), .C(n6990), .Y(n9703) );
  NAND2X1 U2865 ( .A(arr[1401]), .B(n3348), .Y(n6990) );
  OAI21X1 U2866 ( .A(n5507), .B(n3345), .C(n6991), .Y(n9704) );
  NAND2X1 U2867 ( .A(arr[1402]), .B(n3348), .Y(n6991) );
  OAI21X1 U2868 ( .A(n5509), .B(n3346), .C(n6992), .Y(n9705) );
  NAND2X1 U2869 ( .A(arr[1403]), .B(n3348), .Y(n6992) );
  OAI21X1 U2870 ( .A(n5511), .B(n3347), .C(n6993), .Y(n9706) );
  NAND2X1 U2871 ( .A(arr[1404]), .B(n3348), .Y(n6993) );
  OAI21X1 U2872 ( .A(n5513), .B(n3347), .C(n6994), .Y(n9707) );
  NAND2X1 U2873 ( .A(arr[1405]), .B(n3348), .Y(n6994) );
  OAI21X1 U2874 ( .A(n5515), .B(n3347), .C(n6995), .Y(n9708) );
  NAND2X1 U2875 ( .A(arr[1406]), .B(n3348), .Y(n6995) );
  OAI21X1 U2876 ( .A(n5517), .B(n3346), .C(n6996), .Y(n9709) );
  NAND2X1 U2877 ( .A(arr[1407]), .B(n3349), .Y(n6996) );
  OAI21X1 U2878 ( .A(n5519), .B(n3348), .C(n6997), .Y(n9710) );
  NAND2X1 U2879 ( .A(arr[1408]), .B(n3349), .Y(n6997) );
  OAI21X1 U2880 ( .A(n5521), .B(n3348), .C(n6998), .Y(n9711) );
  NAND2X1 U2881 ( .A(arr[1409]), .B(n3349), .Y(n6998) );
  OAI21X1 U2882 ( .A(n5523), .B(n3347), .C(n6999), .Y(n9712) );
  NAND2X1 U2883 ( .A(arr[1410]), .B(n3349), .Y(n6999) );
  OAI21X1 U2884 ( .A(n5525), .B(n3347), .C(n7000), .Y(n9713) );
  NAND2X1 U2885 ( .A(arr[1411]), .B(n3349), .Y(n7000) );
  OAI21X1 U2886 ( .A(n5527), .B(n3347), .C(n7001), .Y(n9714) );
  NAND2X1 U2887 ( .A(arr[1412]), .B(n3349), .Y(n7001) );
  OAI21X1 U2888 ( .A(n5529), .B(n3347), .C(n7002), .Y(n9715) );
  NAND2X1 U2889 ( .A(arr[1413]), .B(n3349), .Y(n7002) );
  OAI21X1 U2890 ( .A(n5531), .B(n3347), .C(n7003), .Y(n9716) );
  NAND2X1 U2891 ( .A(arr[1414]), .B(n3349), .Y(n7003) );
  OAI21X1 U2892 ( .A(n5533), .B(n3347), .C(n7004), .Y(n9717) );
  NAND2X1 U2893 ( .A(arr[1415]), .B(n3349), .Y(n7004) );
  OAI21X1 U2894 ( .A(n5535), .B(n3347), .C(n7005), .Y(n9718) );
  NAND2X1 U2895 ( .A(arr[1416]), .B(n3349), .Y(n7005) );
  OAI21X1 U2896 ( .A(n5537), .B(n3347), .C(n7006), .Y(n9719) );
  NAND2X1 U2897 ( .A(arr[1417]), .B(n3349), .Y(n7006) );
  OAI21X1 U2898 ( .A(n5539), .B(n3347), .C(n7007), .Y(n9720) );
  NAND2X1 U2899 ( .A(arr[1418]), .B(n3349), .Y(n7007) );
  OAI21X1 U2900 ( .A(n5541), .B(n3347), .C(n7008), .Y(n9721) );
  NAND2X1 U2901 ( .A(arr[1419]), .B(n3349), .Y(n7008) );
  OAI21X1 U2902 ( .A(n5543), .B(n3346), .C(n7009), .Y(n9722) );
  NAND2X1 U2903 ( .A(arr[1420]), .B(n3349), .Y(n7009) );
  OAI21X1 U2904 ( .A(n5545), .B(n3346), .C(n7010), .Y(n9723) );
  NAND2X1 U2905 ( .A(arr[1421]), .B(n3349), .Y(n7010) );
  OAI21X1 U2906 ( .A(n5547), .B(n3346), .C(n7011), .Y(n9724) );
  NAND2X1 U2907 ( .A(arr[1422]), .B(n3349), .Y(n7011) );
  OAI21X1 U2908 ( .A(n5549), .B(n3346), .C(n7012), .Y(n9725) );
  NAND2X1 U2909 ( .A(arr[1423]), .B(n3349), .Y(n7012) );
  OAI21X1 U2910 ( .A(n5551), .B(n3346), .C(n7013), .Y(n9726) );
  NAND2X1 U2911 ( .A(arr[1424]), .B(n3350), .Y(n7013) );
  OAI21X1 U2912 ( .A(n5553), .B(n3346), .C(n7014), .Y(n9727) );
  NAND2X1 U2913 ( .A(arr[1425]), .B(n3350), .Y(n7014) );
  OAI21X1 U2914 ( .A(n5555), .B(n3346), .C(n7015), .Y(n9728) );
  NAND2X1 U2915 ( .A(arr[1426]), .B(n3350), .Y(n7015) );
  OAI21X1 U2916 ( .A(n5557), .B(n3346), .C(n7016), .Y(n9729) );
  NAND2X1 U2917 ( .A(arr[1427]), .B(n3350), .Y(n7016) );
  OAI21X1 U2918 ( .A(n5559), .B(n3345), .C(n7017), .Y(n9730) );
  NAND2X1 U2919 ( .A(arr[1428]), .B(n3350), .Y(n7017) );
  OAI21X1 U2920 ( .A(n5561), .B(n3345), .C(n7018), .Y(n9731) );
  NAND2X1 U2921 ( .A(arr[1429]), .B(n3350), .Y(n7018) );
  OAI21X1 U2922 ( .A(n5563), .B(n3345), .C(n7019), .Y(n9732) );
  NAND2X1 U2923 ( .A(arr[1430]), .B(n3350), .Y(n7019) );
  OAI21X1 U2924 ( .A(n5565), .B(n3345), .C(n7020), .Y(n9733) );
  NAND2X1 U2925 ( .A(arr[1431]), .B(n3350), .Y(n7020) );
  OAI21X1 U2926 ( .A(n5567), .B(n3345), .C(n7021), .Y(n9734) );
  NAND2X1 U2927 ( .A(arr[1432]), .B(n3350), .Y(n7021) );
  OAI21X1 U2928 ( .A(n5569), .B(n3345), .C(n7022), .Y(n9735) );
  NAND2X1 U2929 ( .A(arr[1433]), .B(n3348), .Y(n7022) );
  OAI21X1 U2930 ( .A(n5571), .B(n3345), .C(n7023), .Y(n9736) );
  NAND2X1 U2931 ( .A(arr[1434]), .B(n3348), .Y(n7023) );
  NAND2X1 U2932 ( .A(n6939), .B(n5660), .Y(n6982) );
  OAI21X1 U2933 ( .A(n5491), .B(n3339), .C(n7025), .Y(n9737) );
  NAND2X1 U2934 ( .A(arr[1435]), .B(n3342), .Y(n7025) );
  OAI21X1 U2935 ( .A(n5493), .B(n3339), .C(n7026), .Y(n9738) );
  NAND2X1 U2936 ( .A(arr[1436]), .B(n3342), .Y(n7026) );
  OAI21X1 U2937 ( .A(n5495), .B(n3339), .C(n7027), .Y(n9739) );
  NAND2X1 U2938 ( .A(arr[1437]), .B(n3342), .Y(n7027) );
  OAI21X1 U2939 ( .A(n5497), .B(n3339), .C(n7028), .Y(n9740) );
  NAND2X1 U2940 ( .A(arr[1438]), .B(n3342), .Y(n7028) );
  OAI21X1 U2941 ( .A(n5499), .B(n3339), .C(n7029), .Y(n9741) );
  NAND2X1 U2942 ( .A(arr[1439]), .B(n3342), .Y(n7029) );
  OAI21X1 U2943 ( .A(n5501), .B(n3340), .C(n7030), .Y(n9742) );
  NAND2X1 U2944 ( .A(arr[1440]), .B(n3342), .Y(n7030) );
  OAI21X1 U2945 ( .A(n5503), .B(n3340), .C(n7031), .Y(n9743) );
  NAND2X1 U2946 ( .A(arr[1441]), .B(n3342), .Y(n7031) );
  OAI21X1 U2947 ( .A(n5505), .B(n3340), .C(n7032), .Y(n9744) );
  NAND2X1 U2948 ( .A(arr[1442]), .B(n3342), .Y(n7032) );
  OAI21X1 U2949 ( .A(n5507), .B(n3339), .C(n7033), .Y(n9745) );
  NAND2X1 U2950 ( .A(arr[1443]), .B(n3342), .Y(n7033) );
  OAI21X1 U2951 ( .A(n5509), .B(n3340), .C(n7034), .Y(n9746) );
  NAND2X1 U2952 ( .A(arr[1444]), .B(n3342), .Y(n7034) );
  OAI21X1 U2953 ( .A(n5511), .B(n3341), .C(n7035), .Y(n9747) );
  NAND2X1 U2954 ( .A(arr[1445]), .B(n3342), .Y(n7035) );
  OAI21X1 U2955 ( .A(n5513), .B(n3341), .C(n7036), .Y(n9748) );
  NAND2X1 U2956 ( .A(arr[1446]), .B(n3342), .Y(n7036) );
  OAI21X1 U2957 ( .A(n5515), .B(n3341), .C(n7037), .Y(n9749) );
  NAND2X1 U2958 ( .A(arr[1447]), .B(n3342), .Y(n7037) );
  OAI21X1 U2959 ( .A(n5517), .B(n3340), .C(n7038), .Y(n9750) );
  NAND2X1 U2960 ( .A(arr[1448]), .B(n3343), .Y(n7038) );
  OAI21X1 U2961 ( .A(n5519), .B(n3342), .C(n7039), .Y(n9751) );
  NAND2X1 U2962 ( .A(arr[1449]), .B(n3343), .Y(n7039) );
  OAI21X1 U2963 ( .A(n5521), .B(n3342), .C(n7040), .Y(n9752) );
  NAND2X1 U2964 ( .A(arr[1450]), .B(n3343), .Y(n7040) );
  OAI21X1 U2965 ( .A(n5523), .B(n3341), .C(n7041), .Y(n9753) );
  NAND2X1 U2966 ( .A(arr[1451]), .B(n3343), .Y(n7041) );
  OAI21X1 U2967 ( .A(n5525), .B(n3341), .C(n7042), .Y(n9754) );
  NAND2X1 U2968 ( .A(arr[1452]), .B(n3343), .Y(n7042) );
  OAI21X1 U2969 ( .A(n5527), .B(n3341), .C(n7043), .Y(n9755) );
  NAND2X1 U2970 ( .A(arr[1453]), .B(n3343), .Y(n7043) );
  OAI21X1 U2971 ( .A(n5529), .B(n3341), .C(n7044), .Y(n9756) );
  NAND2X1 U2972 ( .A(arr[1454]), .B(n3343), .Y(n7044) );
  OAI21X1 U2973 ( .A(n5531), .B(n3341), .C(n7045), .Y(n9757) );
  NAND2X1 U2974 ( .A(arr[1455]), .B(n3343), .Y(n7045) );
  OAI21X1 U2975 ( .A(n5533), .B(n3341), .C(n7046), .Y(n9758) );
  NAND2X1 U2976 ( .A(arr[1456]), .B(n3343), .Y(n7046) );
  OAI21X1 U2977 ( .A(n5535), .B(n3341), .C(n7047), .Y(n9759) );
  NAND2X1 U2978 ( .A(arr[1457]), .B(n3343), .Y(n7047) );
  OAI21X1 U2979 ( .A(n5537), .B(n3341), .C(n7048), .Y(n9760) );
  NAND2X1 U2980 ( .A(arr[1458]), .B(n3343), .Y(n7048) );
  OAI21X1 U2981 ( .A(n5539), .B(n3341), .C(n7049), .Y(n9761) );
  NAND2X1 U2982 ( .A(arr[1459]), .B(n3343), .Y(n7049) );
  OAI21X1 U2983 ( .A(n5541), .B(n3341), .C(n7050), .Y(n9762) );
  NAND2X1 U2984 ( .A(arr[1460]), .B(n3343), .Y(n7050) );
  OAI21X1 U2985 ( .A(n5543), .B(n3340), .C(n7051), .Y(n9763) );
  NAND2X1 U2986 ( .A(arr[1461]), .B(n3343), .Y(n7051) );
  OAI21X1 U2987 ( .A(n5545), .B(n3340), .C(n7052), .Y(n9764) );
  NAND2X1 U2988 ( .A(arr[1462]), .B(n3343), .Y(n7052) );
  OAI21X1 U2989 ( .A(n5547), .B(n3340), .C(n7053), .Y(n9765) );
  NAND2X1 U2990 ( .A(arr[1463]), .B(n3343), .Y(n7053) );
  OAI21X1 U2991 ( .A(n5549), .B(n3340), .C(n7054), .Y(n9766) );
  NAND2X1 U2992 ( .A(arr[1464]), .B(n3343), .Y(n7054) );
  OAI21X1 U2993 ( .A(n5551), .B(n3340), .C(n7055), .Y(n9767) );
  NAND2X1 U2994 ( .A(arr[1465]), .B(n3344), .Y(n7055) );
  OAI21X1 U2995 ( .A(n5553), .B(n3340), .C(n7056), .Y(n9768) );
  NAND2X1 U2996 ( .A(arr[1466]), .B(n3344), .Y(n7056) );
  OAI21X1 U2997 ( .A(n5555), .B(n3340), .C(n7057), .Y(n9769) );
  NAND2X1 U2998 ( .A(arr[1467]), .B(n3344), .Y(n7057) );
  OAI21X1 U2999 ( .A(n5557), .B(n3340), .C(n7058), .Y(n9770) );
  NAND2X1 U3000 ( .A(arr[1468]), .B(n3344), .Y(n7058) );
  OAI21X1 U3001 ( .A(n5559), .B(n3339), .C(n7059), .Y(n9771) );
  NAND2X1 U3002 ( .A(arr[1469]), .B(n3344), .Y(n7059) );
  OAI21X1 U3003 ( .A(n5561), .B(n3339), .C(n7060), .Y(n9772) );
  NAND2X1 U3004 ( .A(arr[1470]), .B(n3344), .Y(n7060) );
  OAI21X1 U3005 ( .A(n5563), .B(n3339), .C(n7061), .Y(n9773) );
  NAND2X1 U3006 ( .A(arr[1471]), .B(n3344), .Y(n7061) );
  OAI21X1 U3007 ( .A(n5565), .B(n3339), .C(n7062), .Y(n9774) );
  NAND2X1 U3008 ( .A(arr[1472]), .B(n3344), .Y(n7062) );
  OAI21X1 U3009 ( .A(n5567), .B(n3339), .C(n7063), .Y(n9775) );
  NAND2X1 U3010 ( .A(arr[1473]), .B(n3344), .Y(n7063) );
  OAI21X1 U3011 ( .A(n5569), .B(n3339), .C(n7064), .Y(n9776) );
  NAND2X1 U3012 ( .A(arr[1474]), .B(n3342), .Y(n7064) );
  OAI21X1 U3013 ( .A(n5571), .B(n3339), .C(n7065), .Y(n9777) );
  NAND2X1 U3014 ( .A(arr[1475]), .B(n3342), .Y(n7065) );
  NAND2X1 U3015 ( .A(n6939), .B(n5703), .Y(n7024) );
  OAI21X1 U3017 ( .A(n5491), .B(n3333), .C(n7068), .Y(n9778) );
  NAND2X1 U3018 ( .A(arr[1476]), .B(n3336), .Y(n7068) );
  OAI21X1 U3019 ( .A(n5493), .B(n3333), .C(n7069), .Y(n9779) );
  NAND2X1 U3020 ( .A(arr[1477]), .B(n3336), .Y(n7069) );
  OAI21X1 U3021 ( .A(n5495), .B(n3333), .C(n7070), .Y(n9780) );
  NAND2X1 U3022 ( .A(arr[1478]), .B(n3336), .Y(n7070) );
  OAI21X1 U3023 ( .A(n5497), .B(n3333), .C(n7071), .Y(n9781) );
  NAND2X1 U3024 ( .A(arr[1479]), .B(n3336), .Y(n7071) );
  OAI21X1 U3025 ( .A(n5499), .B(n3333), .C(n7072), .Y(n9782) );
  NAND2X1 U3026 ( .A(arr[1480]), .B(n3336), .Y(n7072) );
  OAI21X1 U3027 ( .A(n5501), .B(n3334), .C(n7073), .Y(n9783) );
  NAND2X1 U3028 ( .A(arr[1481]), .B(n3336), .Y(n7073) );
  OAI21X1 U3029 ( .A(n5503), .B(n3334), .C(n7074), .Y(n9784) );
  NAND2X1 U3030 ( .A(arr[1482]), .B(n3336), .Y(n7074) );
  OAI21X1 U3031 ( .A(n5505), .B(n3334), .C(n7075), .Y(n9785) );
  NAND2X1 U3032 ( .A(arr[1483]), .B(n3336), .Y(n7075) );
  OAI21X1 U3033 ( .A(n5507), .B(n3333), .C(n7076), .Y(n9786) );
  NAND2X1 U3034 ( .A(arr[1484]), .B(n3336), .Y(n7076) );
  OAI21X1 U3035 ( .A(n5509), .B(n3334), .C(n7077), .Y(n9787) );
  NAND2X1 U3036 ( .A(arr[1485]), .B(n3336), .Y(n7077) );
  OAI21X1 U3037 ( .A(n5511), .B(n3335), .C(n7078), .Y(n9788) );
  NAND2X1 U3038 ( .A(arr[1486]), .B(n3336), .Y(n7078) );
  OAI21X1 U3039 ( .A(n5513), .B(n3335), .C(n7079), .Y(n9789) );
  NAND2X1 U3040 ( .A(arr[1487]), .B(n3336), .Y(n7079) );
  OAI21X1 U3041 ( .A(n5515), .B(n3335), .C(n7080), .Y(n9790) );
  NAND2X1 U3042 ( .A(arr[1488]), .B(n3336), .Y(n7080) );
  OAI21X1 U3043 ( .A(n5517), .B(n3334), .C(n7081), .Y(n9791) );
  NAND2X1 U3044 ( .A(arr[1489]), .B(n3337), .Y(n7081) );
  OAI21X1 U3045 ( .A(n5519), .B(n3336), .C(n7082), .Y(n9792) );
  NAND2X1 U3046 ( .A(arr[1490]), .B(n3337), .Y(n7082) );
  OAI21X1 U3047 ( .A(n5521), .B(n3336), .C(n7083), .Y(n9793) );
  NAND2X1 U3048 ( .A(arr[1491]), .B(n3337), .Y(n7083) );
  OAI21X1 U3049 ( .A(n5523), .B(n3335), .C(n7084), .Y(n9794) );
  NAND2X1 U3050 ( .A(arr[1492]), .B(n3337), .Y(n7084) );
  OAI21X1 U3051 ( .A(n5525), .B(n3335), .C(n7085), .Y(n9795) );
  NAND2X1 U3052 ( .A(arr[1493]), .B(n3337), .Y(n7085) );
  OAI21X1 U3053 ( .A(n5527), .B(n3335), .C(n7086), .Y(n9796) );
  NAND2X1 U3054 ( .A(arr[1494]), .B(n3337), .Y(n7086) );
  OAI21X1 U3055 ( .A(n5529), .B(n3335), .C(n7087), .Y(n9797) );
  NAND2X1 U3056 ( .A(arr[1495]), .B(n3337), .Y(n7087) );
  OAI21X1 U3057 ( .A(n5531), .B(n3335), .C(n7088), .Y(n9798) );
  NAND2X1 U3058 ( .A(arr[1496]), .B(n3337), .Y(n7088) );
  OAI21X1 U3059 ( .A(n5533), .B(n3335), .C(n7089), .Y(n9799) );
  NAND2X1 U3060 ( .A(arr[1497]), .B(n3337), .Y(n7089) );
  OAI21X1 U3061 ( .A(n5535), .B(n3335), .C(n7090), .Y(n9800) );
  NAND2X1 U3062 ( .A(arr[1498]), .B(n3337), .Y(n7090) );
  OAI21X1 U3063 ( .A(n5537), .B(n3335), .C(n7091), .Y(n9801) );
  NAND2X1 U3064 ( .A(arr[1499]), .B(n3337), .Y(n7091) );
  OAI21X1 U3065 ( .A(n5539), .B(n3335), .C(n7092), .Y(n9802) );
  NAND2X1 U3066 ( .A(arr[1500]), .B(n3337), .Y(n7092) );
  OAI21X1 U3067 ( .A(n5541), .B(n3335), .C(n7093), .Y(n9803) );
  NAND2X1 U3068 ( .A(arr[1501]), .B(n3337), .Y(n7093) );
  OAI21X1 U3069 ( .A(n5543), .B(n3334), .C(n7094), .Y(n9804) );
  NAND2X1 U3070 ( .A(arr[1502]), .B(n3337), .Y(n7094) );
  OAI21X1 U3071 ( .A(n5545), .B(n3334), .C(n7095), .Y(n9805) );
  NAND2X1 U3072 ( .A(arr[1503]), .B(n3337), .Y(n7095) );
  OAI21X1 U3073 ( .A(n5547), .B(n3334), .C(n7096), .Y(n9806) );
  NAND2X1 U3074 ( .A(arr[1504]), .B(n3337), .Y(n7096) );
  OAI21X1 U3075 ( .A(n5549), .B(n3334), .C(n7097), .Y(n9807) );
  NAND2X1 U3076 ( .A(arr[1505]), .B(n3337), .Y(n7097) );
  OAI21X1 U3077 ( .A(n5551), .B(n3334), .C(n7098), .Y(n9808) );
  NAND2X1 U3078 ( .A(arr[1506]), .B(n3338), .Y(n7098) );
  OAI21X1 U3079 ( .A(n5553), .B(n3334), .C(n7099), .Y(n9809) );
  NAND2X1 U3080 ( .A(arr[1507]), .B(n3338), .Y(n7099) );
  OAI21X1 U3081 ( .A(n5555), .B(n3334), .C(n7100), .Y(n9810) );
  NAND2X1 U3082 ( .A(arr[1508]), .B(n3338), .Y(n7100) );
  OAI21X1 U3083 ( .A(n5557), .B(n3334), .C(n7101), .Y(n9811) );
  NAND2X1 U3084 ( .A(arr[1509]), .B(n3338), .Y(n7101) );
  OAI21X1 U3085 ( .A(n5559), .B(n3333), .C(n7102), .Y(n9812) );
  NAND2X1 U3086 ( .A(arr[1510]), .B(n3338), .Y(n7102) );
  OAI21X1 U3087 ( .A(n5561), .B(n3333), .C(n7103), .Y(n9813) );
  NAND2X1 U3088 ( .A(arr[1511]), .B(n3338), .Y(n7103) );
  OAI21X1 U3089 ( .A(n5563), .B(n3333), .C(n7104), .Y(n9814) );
  NAND2X1 U3090 ( .A(arr[1512]), .B(n3338), .Y(n7104) );
  OAI21X1 U3091 ( .A(n5565), .B(n3333), .C(n7105), .Y(n9815) );
  NAND2X1 U3092 ( .A(arr[1513]), .B(n3338), .Y(n7105) );
  OAI21X1 U3093 ( .A(n5567), .B(n3333), .C(n7106), .Y(n9816) );
  NAND2X1 U3094 ( .A(arr[1514]), .B(n3338), .Y(n7106) );
  OAI21X1 U3095 ( .A(n5569), .B(n3333), .C(n7107), .Y(n9817) );
  NAND2X1 U3096 ( .A(arr[1515]), .B(n3336), .Y(n7107) );
  OAI21X1 U3097 ( .A(n5571), .B(n3333), .C(n7108), .Y(n9818) );
  NAND2X1 U3098 ( .A(arr[1516]), .B(n3336), .Y(n7108) );
  NAND2X1 U3099 ( .A(n7109), .B(n5573), .Y(n7067) );
  OAI21X1 U3100 ( .A(n5491), .B(n3327), .C(n7111), .Y(n9819) );
  NAND2X1 U3101 ( .A(arr[1517]), .B(n3330), .Y(n7111) );
  OAI21X1 U3102 ( .A(n5493), .B(n3327), .C(n7112), .Y(n9820) );
  NAND2X1 U3103 ( .A(arr[1518]), .B(n3330), .Y(n7112) );
  OAI21X1 U3104 ( .A(n5495), .B(n3327), .C(n7113), .Y(n9821) );
  NAND2X1 U3105 ( .A(arr[1519]), .B(n3330), .Y(n7113) );
  OAI21X1 U3106 ( .A(n5497), .B(n3327), .C(n7114), .Y(n9822) );
  NAND2X1 U3107 ( .A(arr[1520]), .B(n3330), .Y(n7114) );
  OAI21X1 U3108 ( .A(n5499), .B(n3327), .C(n7115), .Y(n9823) );
  NAND2X1 U3109 ( .A(arr[1521]), .B(n3330), .Y(n7115) );
  OAI21X1 U3110 ( .A(n5501), .B(n3328), .C(n7116), .Y(n9824) );
  NAND2X1 U3111 ( .A(arr[1522]), .B(n3330), .Y(n7116) );
  OAI21X1 U3112 ( .A(n5503), .B(n3328), .C(n7117), .Y(n9825) );
  NAND2X1 U3113 ( .A(arr[1523]), .B(n3330), .Y(n7117) );
  OAI21X1 U3114 ( .A(n5505), .B(n3328), .C(n7118), .Y(n9826) );
  NAND2X1 U3115 ( .A(arr[1524]), .B(n3330), .Y(n7118) );
  OAI21X1 U3116 ( .A(n5507), .B(n3327), .C(n7119), .Y(n9827) );
  NAND2X1 U3117 ( .A(arr[1525]), .B(n3330), .Y(n7119) );
  OAI21X1 U3118 ( .A(n5509), .B(n3328), .C(n7120), .Y(n9828) );
  NAND2X1 U3119 ( .A(arr[1526]), .B(n3330), .Y(n7120) );
  OAI21X1 U3120 ( .A(n5511), .B(n3329), .C(n7121), .Y(n9829) );
  NAND2X1 U3121 ( .A(arr[1527]), .B(n3330), .Y(n7121) );
  OAI21X1 U3122 ( .A(n5513), .B(n3329), .C(n7122), .Y(n9830) );
  NAND2X1 U3123 ( .A(arr[1528]), .B(n3330), .Y(n7122) );
  OAI21X1 U3124 ( .A(n5515), .B(n3329), .C(n7123), .Y(n9831) );
  NAND2X1 U3125 ( .A(arr[1529]), .B(n3330), .Y(n7123) );
  OAI21X1 U3126 ( .A(n5517), .B(n3328), .C(n7124), .Y(n9832) );
  NAND2X1 U3127 ( .A(arr[1530]), .B(n3331), .Y(n7124) );
  OAI21X1 U3128 ( .A(n5519), .B(n3330), .C(n7125), .Y(n9833) );
  NAND2X1 U3129 ( .A(arr[1531]), .B(n3331), .Y(n7125) );
  OAI21X1 U3130 ( .A(n5521), .B(n3330), .C(n7126), .Y(n9834) );
  NAND2X1 U3131 ( .A(arr[1532]), .B(n3331), .Y(n7126) );
  OAI21X1 U3132 ( .A(n5523), .B(n3329), .C(n7127), .Y(n9835) );
  NAND2X1 U3133 ( .A(arr[1533]), .B(n3331), .Y(n7127) );
  OAI21X1 U3134 ( .A(n5525), .B(n3329), .C(n7128), .Y(n9836) );
  NAND2X1 U3135 ( .A(arr[1534]), .B(n3331), .Y(n7128) );
  OAI21X1 U3136 ( .A(n5527), .B(n3329), .C(n7129), .Y(n9837) );
  NAND2X1 U3137 ( .A(arr[1535]), .B(n3331), .Y(n7129) );
  OAI21X1 U3138 ( .A(n5529), .B(n3329), .C(n7130), .Y(n9838) );
  NAND2X1 U3139 ( .A(arr[1536]), .B(n3331), .Y(n7130) );
  OAI21X1 U3140 ( .A(n5531), .B(n3329), .C(n7131), .Y(n9839) );
  NAND2X1 U3141 ( .A(arr[1537]), .B(n3331), .Y(n7131) );
  OAI21X1 U3142 ( .A(n5533), .B(n3329), .C(n7132), .Y(n9840) );
  NAND2X1 U3143 ( .A(arr[1538]), .B(n3331), .Y(n7132) );
  OAI21X1 U3144 ( .A(n5535), .B(n3329), .C(n7133), .Y(n9841) );
  NAND2X1 U3145 ( .A(arr[1539]), .B(n3331), .Y(n7133) );
  OAI21X1 U3146 ( .A(n5537), .B(n3329), .C(n7134), .Y(n9842) );
  NAND2X1 U3147 ( .A(arr[1540]), .B(n3331), .Y(n7134) );
  OAI21X1 U3148 ( .A(n5539), .B(n3329), .C(n7135), .Y(n9843) );
  NAND2X1 U3149 ( .A(arr[1541]), .B(n3331), .Y(n7135) );
  OAI21X1 U3150 ( .A(n5541), .B(n3329), .C(n7136), .Y(n9844) );
  NAND2X1 U3151 ( .A(arr[1542]), .B(n3331), .Y(n7136) );
  OAI21X1 U3152 ( .A(n5543), .B(n3328), .C(n7137), .Y(n9845) );
  NAND2X1 U3153 ( .A(arr[1543]), .B(n3331), .Y(n7137) );
  OAI21X1 U3154 ( .A(n5545), .B(n3328), .C(n7138), .Y(n9846) );
  NAND2X1 U3155 ( .A(arr[1544]), .B(n3331), .Y(n7138) );
  OAI21X1 U3156 ( .A(n5547), .B(n3328), .C(n7139), .Y(n9847) );
  NAND2X1 U3157 ( .A(arr[1545]), .B(n3331), .Y(n7139) );
  OAI21X1 U3158 ( .A(n5549), .B(n3328), .C(n7140), .Y(n9848) );
  NAND2X1 U3159 ( .A(arr[1546]), .B(n3331), .Y(n7140) );
  OAI21X1 U3160 ( .A(n5551), .B(n3328), .C(n7141), .Y(n9849) );
  NAND2X1 U3161 ( .A(arr[1547]), .B(n3332), .Y(n7141) );
  OAI21X1 U3162 ( .A(n5553), .B(n3328), .C(n7142), .Y(n9850) );
  NAND2X1 U3163 ( .A(arr[1548]), .B(n3332), .Y(n7142) );
  OAI21X1 U3164 ( .A(n5555), .B(n3328), .C(n7143), .Y(n9851) );
  NAND2X1 U3165 ( .A(arr[1549]), .B(n3332), .Y(n7143) );
  OAI21X1 U3166 ( .A(n5557), .B(n3328), .C(n7144), .Y(n9852) );
  NAND2X1 U3167 ( .A(arr[1550]), .B(n3332), .Y(n7144) );
  OAI21X1 U3168 ( .A(n5559), .B(n3327), .C(n7145), .Y(n9853) );
  NAND2X1 U3169 ( .A(arr[1551]), .B(n3332), .Y(n7145) );
  OAI21X1 U3170 ( .A(n5561), .B(n3327), .C(n7146), .Y(n9854) );
  NAND2X1 U3171 ( .A(arr[1552]), .B(n3332), .Y(n7146) );
  OAI21X1 U3172 ( .A(n5563), .B(n3327), .C(n7147), .Y(n9855) );
  NAND2X1 U3173 ( .A(arr[1553]), .B(n3332), .Y(n7147) );
  OAI21X1 U3174 ( .A(n5565), .B(n3327), .C(n7148), .Y(n9856) );
  NAND2X1 U3175 ( .A(arr[1554]), .B(n3332), .Y(n7148) );
  OAI21X1 U3176 ( .A(n5567), .B(n3327), .C(n7149), .Y(n9857) );
  NAND2X1 U3177 ( .A(arr[1555]), .B(n3332), .Y(n7149) );
  OAI21X1 U3178 ( .A(n5569), .B(n3327), .C(n7150), .Y(n9858) );
  NAND2X1 U3179 ( .A(arr[1556]), .B(n3330), .Y(n7150) );
  OAI21X1 U3180 ( .A(n5571), .B(n3327), .C(n7151), .Y(n9859) );
  NAND2X1 U3181 ( .A(arr[1557]), .B(n3330), .Y(n7151) );
  NAND2X1 U3182 ( .A(n7109), .B(n5617), .Y(n7110) );
  OAI21X1 U3183 ( .A(n5491), .B(n3321), .C(n7153), .Y(n9860) );
  NAND2X1 U3184 ( .A(arr[1558]), .B(n3324), .Y(n7153) );
  OAI21X1 U3185 ( .A(n5493), .B(n3321), .C(n7154), .Y(n9861) );
  NAND2X1 U3186 ( .A(arr[1559]), .B(n3324), .Y(n7154) );
  OAI21X1 U3187 ( .A(n5495), .B(n3321), .C(n7155), .Y(n9862) );
  NAND2X1 U3188 ( .A(arr[1560]), .B(n3324), .Y(n7155) );
  OAI21X1 U3189 ( .A(n5497), .B(n3321), .C(n7156), .Y(n9863) );
  NAND2X1 U3190 ( .A(arr[1561]), .B(n3324), .Y(n7156) );
  OAI21X1 U3191 ( .A(n5499), .B(n3321), .C(n7157), .Y(n9864) );
  NAND2X1 U3192 ( .A(arr[1562]), .B(n3324), .Y(n7157) );
  OAI21X1 U3193 ( .A(n5501), .B(n3322), .C(n7158), .Y(n9865) );
  NAND2X1 U3194 ( .A(arr[1563]), .B(n3324), .Y(n7158) );
  OAI21X1 U3195 ( .A(n5503), .B(n3322), .C(n7159), .Y(n9866) );
  NAND2X1 U3196 ( .A(arr[1564]), .B(n3324), .Y(n7159) );
  OAI21X1 U3197 ( .A(n5505), .B(n3322), .C(n7160), .Y(n9867) );
  NAND2X1 U3198 ( .A(arr[1565]), .B(n3324), .Y(n7160) );
  OAI21X1 U3199 ( .A(n5507), .B(n3321), .C(n7161), .Y(n9868) );
  NAND2X1 U3200 ( .A(arr[1566]), .B(n3324), .Y(n7161) );
  OAI21X1 U3201 ( .A(n5509), .B(n3322), .C(n7162), .Y(n9869) );
  NAND2X1 U3202 ( .A(arr[1567]), .B(n3324), .Y(n7162) );
  OAI21X1 U3203 ( .A(n5511), .B(n3323), .C(n7163), .Y(n9870) );
  NAND2X1 U3204 ( .A(arr[1568]), .B(n3324), .Y(n7163) );
  OAI21X1 U3205 ( .A(n5513), .B(n3323), .C(n7164), .Y(n9871) );
  NAND2X1 U3206 ( .A(arr[1569]), .B(n3324), .Y(n7164) );
  OAI21X1 U3207 ( .A(n5515), .B(n3323), .C(n7165), .Y(n9872) );
  NAND2X1 U3208 ( .A(arr[1570]), .B(n3324), .Y(n7165) );
  OAI21X1 U3209 ( .A(n5517), .B(n3322), .C(n7166), .Y(n9873) );
  NAND2X1 U3210 ( .A(arr[1571]), .B(n3325), .Y(n7166) );
  OAI21X1 U3211 ( .A(n5519), .B(n3324), .C(n7167), .Y(n9874) );
  NAND2X1 U3212 ( .A(arr[1572]), .B(n3325), .Y(n7167) );
  OAI21X1 U3213 ( .A(n5521), .B(n3324), .C(n7168), .Y(n9875) );
  NAND2X1 U3214 ( .A(arr[1573]), .B(n3325), .Y(n7168) );
  OAI21X1 U3215 ( .A(n5523), .B(n3323), .C(n7169), .Y(n9876) );
  NAND2X1 U3216 ( .A(arr[1574]), .B(n3325), .Y(n7169) );
  OAI21X1 U3217 ( .A(n5525), .B(n3323), .C(n7170), .Y(n9877) );
  NAND2X1 U3218 ( .A(arr[1575]), .B(n3325), .Y(n7170) );
  OAI21X1 U3219 ( .A(n5527), .B(n3323), .C(n7171), .Y(n9878) );
  NAND2X1 U3220 ( .A(arr[1576]), .B(n3325), .Y(n7171) );
  OAI21X1 U3221 ( .A(n5529), .B(n3323), .C(n7172), .Y(n9879) );
  NAND2X1 U3222 ( .A(arr[1577]), .B(n3325), .Y(n7172) );
  OAI21X1 U3223 ( .A(n5531), .B(n3323), .C(n7173), .Y(n9880) );
  NAND2X1 U3224 ( .A(arr[1578]), .B(n3325), .Y(n7173) );
  OAI21X1 U3225 ( .A(n5533), .B(n3323), .C(n7174), .Y(n9881) );
  NAND2X1 U3226 ( .A(arr[1579]), .B(n3325), .Y(n7174) );
  OAI21X1 U3227 ( .A(n5535), .B(n3323), .C(n7175), .Y(n9882) );
  NAND2X1 U3228 ( .A(arr[1580]), .B(n3325), .Y(n7175) );
  OAI21X1 U3229 ( .A(n5537), .B(n3323), .C(n7176), .Y(n9883) );
  NAND2X1 U3230 ( .A(arr[1581]), .B(n3325), .Y(n7176) );
  OAI21X1 U3231 ( .A(n5539), .B(n3323), .C(n7177), .Y(n9884) );
  NAND2X1 U3232 ( .A(arr[1582]), .B(n3325), .Y(n7177) );
  OAI21X1 U3233 ( .A(n5541), .B(n3323), .C(n7178), .Y(n9885) );
  NAND2X1 U3234 ( .A(arr[1583]), .B(n3325), .Y(n7178) );
  OAI21X1 U3235 ( .A(n5543), .B(n3322), .C(n7179), .Y(n9886) );
  NAND2X1 U3236 ( .A(arr[1584]), .B(n3325), .Y(n7179) );
  OAI21X1 U3237 ( .A(n5545), .B(n3322), .C(n7180), .Y(n9887) );
  NAND2X1 U3238 ( .A(arr[1585]), .B(n3325), .Y(n7180) );
  OAI21X1 U3239 ( .A(n5547), .B(n3322), .C(n7181), .Y(n9888) );
  NAND2X1 U3240 ( .A(arr[1586]), .B(n3325), .Y(n7181) );
  OAI21X1 U3241 ( .A(n5549), .B(n3322), .C(n7182), .Y(n9889) );
  NAND2X1 U3242 ( .A(arr[1587]), .B(n3325), .Y(n7182) );
  OAI21X1 U3243 ( .A(n5551), .B(n3322), .C(n7183), .Y(n9890) );
  NAND2X1 U3244 ( .A(arr[1588]), .B(n3326), .Y(n7183) );
  OAI21X1 U3245 ( .A(n5553), .B(n3322), .C(n7184), .Y(n9891) );
  NAND2X1 U3246 ( .A(arr[1589]), .B(n3326), .Y(n7184) );
  OAI21X1 U3247 ( .A(n5555), .B(n3322), .C(n7185), .Y(n9892) );
  NAND2X1 U3248 ( .A(arr[1590]), .B(n3326), .Y(n7185) );
  OAI21X1 U3249 ( .A(n5557), .B(n3322), .C(n7186), .Y(n9893) );
  NAND2X1 U3250 ( .A(arr[1591]), .B(n3326), .Y(n7186) );
  OAI21X1 U3251 ( .A(n5559), .B(n3321), .C(n7187), .Y(n9894) );
  NAND2X1 U3252 ( .A(arr[1592]), .B(n3326), .Y(n7187) );
  OAI21X1 U3253 ( .A(n5561), .B(n3321), .C(n7188), .Y(n9895) );
  NAND2X1 U3254 ( .A(arr[1593]), .B(n3326), .Y(n7188) );
  OAI21X1 U3255 ( .A(n5563), .B(n3321), .C(n7189), .Y(n9896) );
  NAND2X1 U3256 ( .A(arr[1594]), .B(n3326), .Y(n7189) );
  OAI21X1 U3257 ( .A(n5565), .B(n3321), .C(n7190), .Y(n9897) );
  NAND2X1 U3258 ( .A(arr[1595]), .B(n3326), .Y(n7190) );
  OAI21X1 U3259 ( .A(n5567), .B(n3321), .C(n7191), .Y(n9898) );
  NAND2X1 U3260 ( .A(arr[1596]), .B(n3326), .Y(n7191) );
  OAI21X1 U3261 ( .A(n5569), .B(n3321), .C(n7192), .Y(n9899) );
  NAND2X1 U3262 ( .A(arr[1597]), .B(n3324), .Y(n7192) );
  OAI21X1 U3263 ( .A(n5571), .B(n3321), .C(n7193), .Y(n9900) );
  NAND2X1 U3264 ( .A(arr[1598]), .B(n3324), .Y(n7193) );
  NAND2X1 U3265 ( .A(n7109), .B(n5660), .Y(n7152) );
  OAI21X1 U3266 ( .A(n5491), .B(n3315), .C(n7195), .Y(n9901) );
  NAND2X1 U3267 ( .A(arr[1599]), .B(n3318), .Y(n7195) );
  OAI21X1 U3268 ( .A(n5493), .B(n3315), .C(n7196), .Y(n9902) );
  NAND2X1 U3269 ( .A(arr[1600]), .B(n3318), .Y(n7196) );
  OAI21X1 U3270 ( .A(n5495), .B(n3315), .C(n7197), .Y(n9903) );
  NAND2X1 U3271 ( .A(arr[1601]), .B(n3318), .Y(n7197) );
  OAI21X1 U3272 ( .A(n5497), .B(n3315), .C(n7198), .Y(n9904) );
  NAND2X1 U3273 ( .A(arr[1602]), .B(n3318), .Y(n7198) );
  OAI21X1 U3274 ( .A(n5499), .B(n3315), .C(n7199), .Y(n9905) );
  NAND2X1 U3275 ( .A(arr[1603]), .B(n3318), .Y(n7199) );
  OAI21X1 U3276 ( .A(n5501), .B(n3316), .C(n7200), .Y(n9906) );
  NAND2X1 U3277 ( .A(arr[1604]), .B(n3318), .Y(n7200) );
  OAI21X1 U3278 ( .A(n5503), .B(n3316), .C(n7201), .Y(n9907) );
  NAND2X1 U3279 ( .A(arr[1605]), .B(n3318), .Y(n7201) );
  OAI21X1 U3280 ( .A(n5505), .B(n3316), .C(n7202), .Y(n9908) );
  NAND2X1 U3281 ( .A(arr[1606]), .B(n3318), .Y(n7202) );
  OAI21X1 U3282 ( .A(n5507), .B(n3315), .C(n7203), .Y(n9909) );
  NAND2X1 U3283 ( .A(arr[1607]), .B(n3318), .Y(n7203) );
  OAI21X1 U3284 ( .A(n5509), .B(n3316), .C(n7204), .Y(n9910) );
  NAND2X1 U3285 ( .A(arr[1608]), .B(n3318), .Y(n7204) );
  OAI21X1 U3286 ( .A(n5511), .B(n3317), .C(n7205), .Y(n9911) );
  NAND2X1 U3287 ( .A(arr[1609]), .B(n3318), .Y(n7205) );
  OAI21X1 U3288 ( .A(n5513), .B(n3317), .C(n7206), .Y(n9912) );
  NAND2X1 U3289 ( .A(arr[1610]), .B(n3318), .Y(n7206) );
  OAI21X1 U3290 ( .A(n5515), .B(n3317), .C(n7207), .Y(n9913) );
  NAND2X1 U3291 ( .A(arr[1611]), .B(n3318), .Y(n7207) );
  OAI21X1 U3292 ( .A(n5517), .B(n3316), .C(n7208), .Y(n9914) );
  NAND2X1 U3293 ( .A(arr[1612]), .B(n3319), .Y(n7208) );
  OAI21X1 U3294 ( .A(n5519), .B(n3318), .C(n7209), .Y(n9915) );
  NAND2X1 U3295 ( .A(arr[1613]), .B(n3319), .Y(n7209) );
  OAI21X1 U3296 ( .A(n5521), .B(n3318), .C(n7210), .Y(n9916) );
  NAND2X1 U3297 ( .A(arr[1614]), .B(n3319), .Y(n7210) );
  OAI21X1 U3298 ( .A(n5523), .B(n3317), .C(n7211), .Y(n9917) );
  NAND2X1 U3299 ( .A(arr[1615]), .B(n3319), .Y(n7211) );
  OAI21X1 U3300 ( .A(n5525), .B(n3317), .C(n7212), .Y(n9918) );
  NAND2X1 U3301 ( .A(arr[1616]), .B(n3319), .Y(n7212) );
  OAI21X1 U3302 ( .A(n5527), .B(n3317), .C(n7213), .Y(n9919) );
  NAND2X1 U3303 ( .A(arr[1617]), .B(n3319), .Y(n7213) );
  OAI21X1 U3304 ( .A(n5529), .B(n3317), .C(n7214), .Y(n9920) );
  NAND2X1 U3305 ( .A(arr[1618]), .B(n3319), .Y(n7214) );
  OAI21X1 U3306 ( .A(n5531), .B(n3317), .C(n7215), .Y(n9921) );
  NAND2X1 U3307 ( .A(arr[1619]), .B(n3319), .Y(n7215) );
  OAI21X1 U3308 ( .A(n5533), .B(n3317), .C(n7216), .Y(n9922) );
  NAND2X1 U3309 ( .A(arr[1620]), .B(n3319), .Y(n7216) );
  OAI21X1 U3310 ( .A(n5535), .B(n3317), .C(n7217), .Y(n9923) );
  NAND2X1 U3311 ( .A(arr[1621]), .B(n3319), .Y(n7217) );
  OAI21X1 U3312 ( .A(n5537), .B(n3317), .C(n7218), .Y(n9924) );
  NAND2X1 U3313 ( .A(arr[1622]), .B(n3319), .Y(n7218) );
  OAI21X1 U3314 ( .A(n5539), .B(n3317), .C(n7219), .Y(n9925) );
  NAND2X1 U3315 ( .A(arr[1623]), .B(n3319), .Y(n7219) );
  OAI21X1 U3316 ( .A(n5541), .B(n3317), .C(n7220), .Y(n9926) );
  NAND2X1 U3317 ( .A(arr[1624]), .B(n3319), .Y(n7220) );
  OAI21X1 U3318 ( .A(n5543), .B(n3316), .C(n7221), .Y(n9927) );
  NAND2X1 U3319 ( .A(arr[1625]), .B(n3319), .Y(n7221) );
  OAI21X1 U3320 ( .A(n5545), .B(n3316), .C(n7222), .Y(n9928) );
  NAND2X1 U3321 ( .A(arr[1626]), .B(n3319), .Y(n7222) );
  OAI21X1 U3322 ( .A(n5547), .B(n3316), .C(n7223), .Y(n9929) );
  NAND2X1 U3323 ( .A(arr[1627]), .B(n3319), .Y(n7223) );
  OAI21X1 U3324 ( .A(n5549), .B(n3316), .C(n7224), .Y(n9930) );
  NAND2X1 U3325 ( .A(arr[1628]), .B(n3319), .Y(n7224) );
  OAI21X1 U3326 ( .A(n5551), .B(n3316), .C(n7225), .Y(n9931) );
  NAND2X1 U3327 ( .A(arr[1629]), .B(n3320), .Y(n7225) );
  OAI21X1 U3328 ( .A(n5553), .B(n3316), .C(n7226), .Y(n9932) );
  NAND2X1 U3329 ( .A(arr[1630]), .B(n3320), .Y(n7226) );
  OAI21X1 U3330 ( .A(n5555), .B(n3316), .C(n7227), .Y(n9933) );
  NAND2X1 U3331 ( .A(arr[1631]), .B(n3320), .Y(n7227) );
  OAI21X1 U3332 ( .A(n5557), .B(n3316), .C(n7228), .Y(n9934) );
  NAND2X1 U3333 ( .A(arr[1632]), .B(n3320), .Y(n7228) );
  OAI21X1 U3334 ( .A(n5559), .B(n3315), .C(n7229), .Y(n9935) );
  NAND2X1 U3335 ( .A(arr[1633]), .B(n3320), .Y(n7229) );
  OAI21X1 U3336 ( .A(n5561), .B(n3315), .C(n7230), .Y(n9936) );
  NAND2X1 U3337 ( .A(arr[1634]), .B(n3320), .Y(n7230) );
  OAI21X1 U3338 ( .A(n5563), .B(n3315), .C(n7231), .Y(n9937) );
  NAND2X1 U3339 ( .A(arr[1635]), .B(n3320), .Y(n7231) );
  OAI21X1 U3340 ( .A(n5565), .B(n3315), .C(n7232), .Y(n9938) );
  NAND2X1 U3341 ( .A(arr[1636]), .B(n3320), .Y(n7232) );
  OAI21X1 U3342 ( .A(n5567), .B(n3315), .C(n7233), .Y(n9939) );
  NAND2X1 U3343 ( .A(arr[1637]), .B(n3320), .Y(n7233) );
  OAI21X1 U3344 ( .A(n5569), .B(n3315), .C(n7234), .Y(n9940) );
  NAND2X1 U3345 ( .A(arr[1638]), .B(n3318), .Y(n7234) );
  OAI21X1 U3346 ( .A(n5571), .B(n3315), .C(n7235), .Y(n9941) );
  NAND2X1 U3347 ( .A(arr[1639]), .B(n3318), .Y(n7235) );
  NAND2X1 U3348 ( .A(n7109), .B(n5703), .Y(n7194) );
  OAI21X1 U3350 ( .A(n5491), .B(n3309), .C(n7237), .Y(n9942) );
  NAND2X1 U3351 ( .A(arr[1640]), .B(n3312), .Y(n7237) );
  OAI21X1 U3352 ( .A(n5493), .B(n3309), .C(n7238), .Y(n9943) );
  NAND2X1 U3353 ( .A(arr[1641]), .B(n3312), .Y(n7238) );
  OAI21X1 U3354 ( .A(n5495), .B(n3309), .C(n7239), .Y(n9944) );
  NAND2X1 U3355 ( .A(arr[1642]), .B(n3312), .Y(n7239) );
  OAI21X1 U3356 ( .A(n5497), .B(n3309), .C(n7240), .Y(n9945) );
  NAND2X1 U3357 ( .A(arr[1643]), .B(n3312), .Y(n7240) );
  OAI21X1 U3358 ( .A(n5499), .B(n3309), .C(n7241), .Y(n9946) );
  NAND2X1 U3359 ( .A(arr[1644]), .B(n3312), .Y(n7241) );
  OAI21X1 U3360 ( .A(n5501), .B(n3310), .C(n7242), .Y(n9947) );
  NAND2X1 U3361 ( .A(arr[1645]), .B(n3312), .Y(n7242) );
  OAI21X1 U3362 ( .A(n5503), .B(n3310), .C(n7243), .Y(n9948) );
  NAND2X1 U3363 ( .A(arr[1646]), .B(n3312), .Y(n7243) );
  OAI21X1 U3364 ( .A(n5505), .B(n3310), .C(n7244), .Y(n9949) );
  NAND2X1 U3365 ( .A(arr[1647]), .B(n3312), .Y(n7244) );
  OAI21X1 U3366 ( .A(n5507), .B(n3309), .C(n7245), .Y(n9950) );
  NAND2X1 U3367 ( .A(arr[1648]), .B(n3312), .Y(n7245) );
  OAI21X1 U3368 ( .A(n5509), .B(n3310), .C(n7246), .Y(n9951) );
  NAND2X1 U3369 ( .A(arr[1649]), .B(n3312), .Y(n7246) );
  OAI21X1 U3370 ( .A(n5511), .B(n3311), .C(n7247), .Y(n9952) );
  NAND2X1 U3371 ( .A(arr[1650]), .B(n3312), .Y(n7247) );
  OAI21X1 U3372 ( .A(n5513), .B(n3311), .C(n7248), .Y(n9953) );
  NAND2X1 U3373 ( .A(arr[1651]), .B(n3312), .Y(n7248) );
  OAI21X1 U3374 ( .A(n5515), .B(n3311), .C(n7249), .Y(n9954) );
  NAND2X1 U3375 ( .A(arr[1652]), .B(n3312), .Y(n7249) );
  OAI21X1 U3376 ( .A(n5517), .B(n3310), .C(n7250), .Y(n9955) );
  NAND2X1 U3377 ( .A(arr[1653]), .B(n3313), .Y(n7250) );
  OAI21X1 U3378 ( .A(n5519), .B(n3312), .C(n7251), .Y(n9956) );
  NAND2X1 U3379 ( .A(arr[1654]), .B(n3313), .Y(n7251) );
  OAI21X1 U3380 ( .A(n5521), .B(n3312), .C(n7252), .Y(n9957) );
  NAND2X1 U3381 ( .A(arr[1655]), .B(n3313), .Y(n7252) );
  OAI21X1 U3382 ( .A(n5523), .B(n3311), .C(n7253), .Y(n9958) );
  NAND2X1 U3383 ( .A(arr[1656]), .B(n3313), .Y(n7253) );
  OAI21X1 U3384 ( .A(n5525), .B(n3311), .C(n7254), .Y(n9959) );
  NAND2X1 U3385 ( .A(arr[1657]), .B(n3313), .Y(n7254) );
  OAI21X1 U3386 ( .A(n5527), .B(n3311), .C(n7255), .Y(n9960) );
  NAND2X1 U3387 ( .A(arr[1658]), .B(n3313), .Y(n7255) );
  OAI21X1 U3388 ( .A(n5529), .B(n3311), .C(n7256), .Y(n9961) );
  NAND2X1 U3389 ( .A(arr[1659]), .B(n3313), .Y(n7256) );
  OAI21X1 U3390 ( .A(n5531), .B(n3311), .C(n7257), .Y(n9962) );
  NAND2X1 U3391 ( .A(arr[1660]), .B(n3313), .Y(n7257) );
  OAI21X1 U3392 ( .A(n5533), .B(n3311), .C(n7258), .Y(n9963) );
  NAND2X1 U3393 ( .A(arr[1661]), .B(n3313), .Y(n7258) );
  OAI21X1 U3394 ( .A(n5535), .B(n3311), .C(n7259), .Y(n9964) );
  NAND2X1 U3395 ( .A(arr[1662]), .B(n3313), .Y(n7259) );
  OAI21X1 U3396 ( .A(n5537), .B(n3311), .C(n7260), .Y(n9965) );
  NAND2X1 U3397 ( .A(arr[1663]), .B(n3313), .Y(n7260) );
  OAI21X1 U3398 ( .A(n5539), .B(n3311), .C(n7261), .Y(n9966) );
  NAND2X1 U3399 ( .A(arr[1664]), .B(n3313), .Y(n7261) );
  OAI21X1 U3400 ( .A(n5541), .B(n3311), .C(n7262), .Y(n9967) );
  NAND2X1 U3401 ( .A(arr[1665]), .B(n3313), .Y(n7262) );
  OAI21X1 U3402 ( .A(n5543), .B(n3310), .C(n7263), .Y(n9968) );
  NAND2X1 U3403 ( .A(arr[1666]), .B(n3313), .Y(n7263) );
  OAI21X1 U3404 ( .A(n5545), .B(n3310), .C(n7264), .Y(n9969) );
  NAND2X1 U3405 ( .A(arr[1667]), .B(n3313), .Y(n7264) );
  OAI21X1 U3406 ( .A(n5547), .B(n3310), .C(n7265), .Y(n9970) );
  NAND2X1 U3407 ( .A(arr[1668]), .B(n3313), .Y(n7265) );
  OAI21X1 U3408 ( .A(n5549), .B(n3310), .C(n7266), .Y(n9971) );
  NAND2X1 U3409 ( .A(arr[1669]), .B(n3313), .Y(n7266) );
  OAI21X1 U3410 ( .A(n5551), .B(n3310), .C(n7267), .Y(n9972) );
  NAND2X1 U3411 ( .A(arr[1670]), .B(n3314), .Y(n7267) );
  OAI21X1 U3412 ( .A(n5553), .B(n3310), .C(n7268), .Y(n9973) );
  NAND2X1 U3413 ( .A(arr[1671]), .B(n3314), .Y(n7268) );
  OAI21X1 U3414 ( .A(n5555), .B(n3310), .C(n7269), .Y(n9974) );
  NAND2X1 U3415 ( .A(arr[1672]), .B(n3314), .Y(n7269) );
  OAI21X1 U3416 ( .A(n5557), .B(n3310), .C(n7270), .Y(n9975) );
  NAND2X1 U3417 ( .A(arr[1673]), .B(n3314), .Y(n7270) );
  OAI21X1 U3418 ( .A(n5559), .B(n3309), .C(n7271), .Y(n9976) );
  NAND2X1 U3419 ( .A(arr[1674]), .B(n3314), .Y(n7271) );
  OAI21X1 U3420 ( .A(n5561), .B(n3309), .C(n7272), .Y(n9977) );
  NAND2X1 U3421 ( .A(arr[1675]), .B(n3314), .Y(n7272) );
  OAI21X1 U3422 ( .A(n5563), .B(n3309), .C(n7273), .Y(n9978) );
  NAND2X1 U3423 ( .A(arr[1676]), .B(n3314), .Y(n7273) );
  OAI21X1 U3424 ( .A(n5565), .B(n3309), .C(n7274), .Y(n9979) );
  NAND2X1 U3425 ( .A(arr[1677]), .B(n3314), .Y(n7274) );
  OAI21X1 U3426 ( .A(n5567), .B(n3309), .C(n7275), .Y(n9980) );
  NAND2X1 U3427 ( .A(arr[1678]), .B(n3314), .Y(n7275) );
  OAI21X1 U3428 ( .A(n5569), .B(n3309), .C(n7276), .Y(n9981) );
  NAND2X1 U3429 ( .A(arr[1679]), .B(n3312), .Y(n7276) );
  OAI21X1 U3430 ( .A(n5571), .B(n3309), .C(n7277), .Y(n9982) );
  NAND2X1 U3431 ( .A(arr[1680]), .B(n3312), .Y(n7277) );
  NAND2X1 U3432 ( .A(n7278), .B(n5573), .Y(n7236) );
  OAI21X1 U3433 ( .A(n5491), .B(n3303), .C(n7280), .Y(n9983) );
  NAND2X1 U3434 ( .A(arr[1681]), .B(n3306), .Y(n7280) );
  OAI21X1 U3435 ( .A(n5493), .B(n3303), .C(n7281), .Y(n9984) );
  NAND2X1 U3436 ( .A(arr[1682]), .B(n3306), .Y(n7281) );
  OAI21X1 U3437 ( .A(n5495), .B(n3303), .C(n7282), .Y(n9985) );
  NAND2X1 U3438 ( .A(arr[1683]), .B(n3306), .Y(n7282) );
  OAI21X1 U3439 ( .A(n5497), .B(n3303), .C(n7283), .Y(n9986) );
  NAND2X1 U3440 ( .A(arr[1684]), .B(n3306), .Y(n7283) );
  OAI21X1 U3441 ( .A(n5499), .B(n3303), .C(n7284), .Y(n9987) );
  NAND2X1 U3442 ( .A(arr[1685]), .B(n3306), .Y(n7284) );
  OAI21X1 U3443 ( .A(n5501), .B(n3304), .C(n7285), .Y(n9988) );
  NAND2X1 U3444 ( .A(arr[1686]), .B(n3306), .Y(n7285) );
  OAI21X1 U3445 ( .A(n5503), .B(n3304), .C(n7286), .Y(n9989) );
  NAND2X1 U3446 ( .A(arr[1687]), .B(n3306), .Y(n7286) );
  OAI21X1 U3447 ( .A(n5505), .B(n3304), .C(n7287), .Y(n9990) );
  NAND2X1 U3448 ( .A(arr[1688]), .B(n3306), .Y(n7287) );
  OAI21X1 U3449 ( .A(n5507), .B(n3303), .C(n7288), .Y(n9991) );
  NAND2X1 U3450 ( .A(arr[1689]), .B(n3306), .Y(n7288) );
  OAI21X1 U3451 ( .A(n5509), .B(n3304), .C(n7289), .Y(n9992) );
  NAND2X1 U3452 ( .A(arr[1690]), .B(n3306), .Y(n7289) );
  OAI21X1 U3453 ( .A(n5511), .B(n3305), .C(n7290), .Y(n9993) );
  NAND2X1 U3454 ( .A(arr[1691]), .B(n3306), .Y(n7290) );
  OAI21X1 U3455 ( .A(n5513), .B(n3305), .C(n7291), .Y(n9994) );
  NAND2X1 U3456 ( .A(arr[1692]), .B(n3306), .Y(n7291) );
  OAI21X1 U3457 ( .A(n5515), .B(n3305), .C(n7292), .Y(n9995) );
  NAND2X1 U3458 ( .A(arr[1693]), .B(n3306), .Y(n7292) );
  OAI21X1 U3459 ( .A(n5517), .B(n3304), .C(n7293), .Y(n9996) );
  NAND2X1 U3460 ( .A(arr[1694]), .B(n3307), .Y(n7293) );
  OAI21X1 U3461 ( .A(n5519), .B(n3306), .C(n7294), .Y(n9997) );
  NAND2X1 U3462 ( .A(arr[1695]), .B(n3307), .Y(n7294) );
  OAI21X1 U3463 ( .A(n5521), .B(n3306), .C(n7295), .Y(n9998) );
  NAND2X1 U3464 ( .A(arr[1696]), .B(n3307), .Y(n7295) );
  OAI21X1 U3465 ( .A(n5523), .B(n3305), .C(n7296), .Y(n9999) );
  NAND2X1 U3466 ( .A(arr[1697]), .B(n3307), .Y(n7296) );
  OAI21X1 U3467 ( .A(n5525), .B(n3305), .C(n7297), .Y(n10000) );
  NAND2X1 U3468 ( .A(arr[1698]), .B(n3307), .Y(n7297) );
  OAI21X1 U3469 ( .A(n5527), .B(n3305), .C(n7298), .Y(n10001) );
  NAND2X1 U3470 ( .A(arr[1699]), .B(n3307), .Y(n7298) );
  OAI21X1 U3471 ( .A(n5529), .B(n3305), .C(n7299), .Y(n10002) );
  NAND2X1 U3472 ( .A(arr[1700]), .B(n3307), .Y(n7299) );
  OAI21X1 U3473 ( .A(n5531), .B(n3305), .C(n7300), .Y(n10003) );
  NAND2X1 U3474 ( .A(arr[1701]), .B(n3307), .Y(n7300) );
  OAI21X1 U3475 ( .A(n5533), .B(n3305), .C(n7301), .Y(n10004) );
  NAND2X1 U3476 ( .A(arr[1702]), .B(n3307), .Y(n7301) );
  OAI21X1 U3477 ( .A(n5535), .B(n3305), .C(n7302), .Y(n10005) );
  NAND2X1 U3478 ( .A(arr[1703]), .B(n3307), .Y(n7302) );
  OAI21X1 U3479 ( .A(n5537), .B(n3305), .C(n7303), .Y(n10006) );
  NAND2X1 U3480 ( .A(arr[1704]), .B(n3307), .Y(n7303) );
  OAI21X1 U3481 ( .A(n5539), .B(n3305), .C(n7304), .Y(n10007) );
  NAND2X1 U3482 ( .A(arr[1705]), .B(n3307), .Y(n7304) );
  OAI21X1 U3483 ( .A(n5541), .B(n3305), .C(n7305), .Y(n10008) );
  NAND2X1 U3484 ( .A(arr[1706]), .B(n3307), .Y(n7305) );
  OAI21X1 U3485 ( .A(n5543), .B(n3304), .C(n7306), .Y(n10009) );
  NAND2X1 U3486 ( .A(arr[1707]), .B(n3307), .Y(n7306) );
  OAI21X1 U3487 ( .A(n5545), .B(n3304), .C(n7307), .Y(n10010) );
  NAND2X1 U3488 ( .A(arr[1708]), .B(n3307), .Y(n7307) );
  OAI21X1 U3489 ( .A(n5547), .B(n3304), .C(n7308), .Y(n10011) );
  NAND2X1 U3490 ( .A(arr[1709]), .B(n3307), .Y(n7308) );
  OAI21X1 U3491 ( .A(n5549), .B(n3304), .C(n7309), .Y(n10012) );
  NAND2X1 U3492 ( .A(arr[1710]), .B(n3307), .Y(n7309) );
  OAI21X1 U3493 ( .A(n5551), .B(n3304), .C(n7310), .Y(n10013) );
  NAND2X1 U3494 ( .A(arr[1711]), .B(n3308), .Y(n7310) );
  OAI21X1 U3495 ( .A(n5553), .B(n3304), .C(n7311), .Y(n10014) );
  NAND2X1 U3496 ( .A(arr[1712]), .B(n3308), .Y(n7311) );
  OAI21X1 U3497 ( .A(n5555), .B(n3304), .C(n7312), .Y(n10015) );
  NAND2X1 U3498 ( .A(arr[1713]), .B(n3308), .Y(n7312) );
  OAI21X1 U3499 ( .A(n5557), .B(n3304), .C(n7313), .Y(n10016) );
  NAND2X1 U3500 ( .A(arr[1714]), .B(n3308), .Y(n7313) );
  OAI21X1 U3501 ( .A(n5559), .B(n3303), .C(n7314), .Y(n10017) );
  NAND2X1 U3502 ( .A(arr[1715]), .B(n3308), .Y(n7314) );
  OAI21X1 U3503 ( .A(n5561), .B(n3303), .C(n7315), .Y(n10018) );
  NAND2X1 U3504 ( .A(arr[1716]), .B(n3308), .Y(n7315) );
  OAI21X1 U3505 ( .A(n5563), .B(n3303), .C(n7316), .Y(n10019) );
  NAND2X1 U3506 ( .A(arr[1717]), .B(n3308), .Y(n7316) );
  OAI21X1 U3507 ( .A(n5565), .B(n3303), .C(n7317), .Y(n10020) );
  NAND2X1 U3508 ( .A(arr[1718]), .B(n3308), .Y(n7317) );
  OAI21X1 U3509 ( .A(n5567), .B(n3303), .C(n7318), .Y(n10021) );
  NAND2X1 U3510 ( .A(arr[1719]), .B(n3308), .Y(n7318) );
  OAI21X1 U3511 ( .A(n5569), .B(n3303), .C(n7319), .Y(n10022) );
  NAND2X1 U3512 ( .A(arr[1720]), .B(n3306), .Y(n7319) );
  OAI21X1 U3513 ( .A(n5571), .B(n3303), .C(n7320), .Y(n10023) );
  NAND2X1 U3514 ( .A(arr[1721]), .B(n3306), .Y(n7320) );
  NAND2X1 U3515 ( .A(n7278), .B(n5617), .Y(n7279) );
  OAI21X1 U3516 ( .A(n5491), .B(n3297), .C(n7322), .Y(n10024) );
  NAND2X1 U3517 ( .A(arr[1722]), .B(n3300), .Y(n7322) );
  OAI21X1 U3518 ( .A(n5493), .B(n3297), .C(n7323), .Y(n10025) );
  NAND2X1 U3519 ( .A(arr[1723]), .B(n3300), .Y(n7323) );
  OAI21X1 U3520 ( .A(n5495), .B(n3297), .C(n7324), .Y(n10026) );
  NAND2X1 U3521 ( .A(arr[1724]), .B(n3300), .Y(n7324) );
  OAI21X1 U3522 ( .A(n5497), .B(n3297), .C(n7325), .Y(n10027) );
  NAND2X1 U3523 ( .A(arr[1725]), .B(n3300), .Y(n7325) );
  OAI21X1 U3524 ( .A(n5499), .B(n3297), .C(n7326), .Y(n10028) );
  NAND2X1 U3525 ( .A(arr[1726]), .B(n3300), .Y(n7326) );
  OAI21X1 U3526 ( .A(n5501), .B(n3298), .C(n7327), .Y(n10029) );
  NAND2X1 U3527 ( .A(arr[1727]), .B(n3300), .Y(n7327) );
  OAI21X1 U3528 ( .A(n5503), .B(n3298), .C(n7328), .Y(n10030) );
  NAND2X1 U3529 ( .A(arr[1728]), .B(n3300), .Y(n7328) );
  OAI21X1 U3530 ( .A(n5505), .B(n3298), .C(n7329), .Y(n10031) );
  NAND2X1 U3531 ( .A(arr[1729]), .B(n3300), .Y(n7329) );
  OAI21X1 U3532 ( .A(n5507), .B(n3297), .C(n7330), .Y(n10032) );
  NAND2X1 U3533 ( .A(arr[1730]), .B(n3300), .Y(n7330) );
  OAI21X1 U3534 ( .A(n5509), .B(n3298), .C(n7331), .Y(n10033) );
  NAND2X1 U3535 ( .A(arr[1731]), .B(n3300), .Y(n7331) );
  OAI21X1 U3536 ( .A(n5511), .B(n3299), .C(n7332), .Y(n10034) );
  NAND2X1 U3537 ( .A(arr[1732]), .B(n3300), .Y(n7332) );
  OAI21X1 U3538 ( .A(n5513), .B(n3299), .C(n7333), .Y(n10035) );
  NAND2X1 U3539 ( .A(arr[1733]), .B(n3300), .Y(n7333) );
  OAI21X1 U3540 ( .A(n5515), .B(n3299), .C(n7334), .Y(n10036) );
  NAND2X1 U3541 ( .A(arr[1734]), .B(n3300), .Y(n7334) );
  OAI21X1 U3542 ( .A(n5517), .B(n3298), .C(n7335), .Y(n10037) );
  NAND2X1 U3543 ( .A(arr[1735]), .B(n3301), .Y(n7335) );
  OAI21X1 U3544 ( .A(n5519), .B(n3300), .C(n7336), .Y(n10038) );
  NAND2X1 U3545 ( .A(arr[1736]), .B(n3301), .Y(n7336) );
  OAI21X1 U3546 ( .A(n5521), .B(n3300), .C(n7337), .Y(n10039) );
  NAND2X1 U3547 ( .A(arr[1737]), .B(n3301), .Y(n7337) );
  OAI21X1 U3548 ( .A(n5523), .B(n3299), .C(n7338), .Y(n10040) );
  NAND2X1 U3549 ( .A(arr[1738]), .B(n3301), .Y(n7338) );
  OAI21X1 U3550 ( .A(n5525), .B(n3299), .C(n7339), .Y(n10041) );
  NAND2X1 U3551 ( .A(arr[1739]), .B(n3301), .Y(n7339) );
  OAI21X1 U3552 ( .A(n5527), .B(n3299), .C(n7340), .Y(n10042) );
  NAND2X1 U3553 ( .A(arr[1740]), .B(n3301), .Y(n7340) );
  OAI21X1 U3554 ( .A(n5529), .B(n3299), .C(n7341), .Y(n10043) );
  NAND2X1 U3555 ( .A(arr[1741]), .B(n3301), .Y(n7341) );
  OAI21X1 U3556 ( .A(n5531), .B(n3299), .C(n7342), .Y(n10044) );
  NAND2X1 U3557 ( .A(arr[1742]), .B(n3301), .Y(n7342) );
  OAI21X1 U3558 ( .A(n5533), .B(n3299), .C(n7343), .Y(n10045) );
  NAND2X1 U3559 ( .A(arr[1743]), .B(n3301), .Y(n7343) );
  OAI21X1 U3560 ( .A(n5535), .B(n3299), .C(n7344), .Y(n10046) );
  NAND2X1 U3561 ( .A(arr[1744]), .B(n3301), .Y(n7344) );
  OAI21X1 U3562 ( .A(n5537), .B(n3299), .C(n7345), .Y(n10047) );
  NAND2X1 U3563 ( .A(arr[1745]), .B(n3301), .Y(n7345) );
  OAI21X1 U3564 ( .A(n5539), .B(n3299), .C(n7346), .Y(n10048) );
  NAND2X1 U3565 ( .A(arr[1746]), .B(n3301), .Y(n7346) );
  OAI21X1 U3566 ( .A(n5541), .B(n3299), .C(n7347), .Y(n10049) );
  NAND2X1 U3567 ( .A(arr[1747]), .B(n3301), .Y(n7347) );
  OAI21X1 U3568 ( .A(n5543), .B(n3298), .C(n7348), .Y(n10050) );
  NAND2X1 U3569 ( .A(arr[1748]), .B(n3301), .Y(n7348) );
  OAI21X1 U3570 ( .A(n5545), .B(n3298), .C(n7349), .Y(n10051) );
  NAND2X1 U3571 ( .A(arr[1749]), .B(n3301), .Y(n7349) );
  OAI21X1 U3572 ( .A(n5547), .B(n3298), .C(n7350), .Y(n10052) );
  NAND2X1 U3573 ( .A(arr[1750]), .B(n3301), .Y(n7350) );
  OAI21X1 U3574 ( .A(n5549), .B(n3298), .C(n7351), .Y(n10053) );
  NAND2X1 U3575 ( .A(arr[1751]), .B(n3301), .Y(n7351) );
  OAI21X1 U3576 ( .A(n5551), .B(n3298), .C(n7352), .Y(n10054) );
  NAND2X1 U3577 ( .A(arr[1752]), .B(n3302), .Y(n7352) );
  OAI21X1 U3578 ( .A(n5553), .B(n3298), .C(n7353), .Y(n10055) );
  NAND2X1 U3579 ( .A(arr[1753]), .B(n3302), .Y(n7353) );
  OAI21X1 U3580 ( .A(n5555), .B(n3298), .C(n7354), .Y(n10056) );
  NAND2X1 U3581 ( .A(arr[1754]), .B(n3302), .Y(n7354) );
  OAI21X1 U3582 ( .A(n5557), .B(n3298), .C(n7355), .Y(n10057) );
  NAND2X1 U3583 ( .A(arr[1755]), .B(n3302), .Y(n7355) );
  OAI21X1 U3584 ( .A(n5559), .B(n3297), .C(n7356), .Y(n10058) );
  NAND2X1 U3585 ( .A(arr[1756]), .B(n3302), .Y(n7356) );
  OAI21X1 U3586 ( .A(n5561), .B(n3297), .C(n7357), .Y(n10059) );
  NAND2X1 U3587 ( .A(arr[1757]), .B(n3302), .Y(n7357) );
  OAI21X1 U3588 ( .A(n5563), .B(n3297), .C(n7358), .Y(n10060) );
  NAND2X1 U3589 ( .A(arr[1758]), .B(n3302), .Y(n7358) );
  OAI21X1 U3590 ( .A(n5565), .B(n3297), .C(n7359), .Y(n10061) );
  NAND2X1 U3591 ( .A(arr[1759]), .B(n3302), .Y(n7359) );
  OAI21X1 U3592 ( .A(n5567), .B(n3297), .C(n7360), .Y(n10062) );
  NAND2X1 U3593 ( .A(arr[1760]), .B(n3302), .Y(n7360) );
  OAI21X1 U3594 ( .A(n5569), .B(n3297), .C(n7361), .Y(n10063) );
  NAND2X1 U3595 ( .A(arr[1761]), .B(n3300), .Y(n7361) );
  OAI21X1 U3596 ( .A(n5571), .B(n3297), .C(n7362), .Y(n10064) );
  NAND2X1 U3597 ( .A(arr[1762]), .B(n3300), .Y(n7362) );
  NAND2X1 U3598 ( .A(n7278), .B(n5660), .Y(n7321) );
  OAI21X1 U3599 ( .A(n5491), .B(n3291), .C(n7364), .Y(n10065) );
  NAND2X1 U3600 ( .A(arr[1763]), .B(n3294), .Y(n7364) );
  OAI21X1 U3601 ( .A(n5493), .B(n3291), .C(n7365), .Y(n10066) );
  NAND2X1 U3602 ( .A(arr[1764]), .B(n3294), .Y(n7365) );
  OAI21X1 U3603 ( .A(n5495), .B(n3291), .C(n7366), .Y(n10067) );
  NAND2X1 U3604 ( .A(arr[1765]), .B(n3294), .Y(n7366) );
  OAI21X1 U3605 ( .A(n5497), .B(n3291), .C(n7367), .Y(n10068) );
  NAND2X1 U3606 ( .A(arr[1766]), .B(n3294), .Y(n7367) );
  OAI21X1 U3607 ( .A(n5499), .B(n3291), .C(n7368), .Y(n10069) );
  NAND2X1 U3608 ( .A(arr[1767]), .B(n3294), .Y(n7368) );
  OAI21X1 U3609 ( .A(n5501), .B(n3292), .C(n7369), .Y(n10070) );
  NAND2X1 U3610 ( .A(arr[1768]), .B(n3294), .Y(n7369) );
  OAI21X1 U3611 ( .A(n5503), .B(n3292), .C(n7370), .Y(n10071) );
  NAND2X1 U3612 ( .A(arr[1769]), .B(n3294), .Y(n7370) );
  OAI21X1 U3613 ( .A(n5505), .B(n3292), .C(n7371), .Y(n10072) );
  NAND2X1 U3614 ( .A(arr[1770]), .B(n3294), .Y(n7371) );
  OAI21X1 U3615 ( .A(n5507), .B(n3291), .C(n7372), .Y(n10073) );
  NAND2X1 U3616 ( .A(arr[1771]), .B(n3294), .Y(n7372) );
  OAI21X1 U3617 ( .A(n5509), .B(n3292), .C(n7373), .Y(n10074) );
  NAND2X1 U3618 ( .A(arr[1772]), .B(n3294), .Y(n7373) );
  OAI21X1 U3619 ( .A(n5511), .B(n3293), .C(n7374), .Y(n10075) );
  NAND2X1 U3620 ( .A(arr[1773]), .B(n3294), .Y(n7374) );
  OAI21X1 U3621 ( .A(n5513), .B(n3293), .C(n7375), .Y(n10076) );
  NAND2X1 U3622 ( .A(arr[1774]), .B(n3294), .Y(n7375) );
  OAI21X1 U3623 ( .A(n5515), .B(n3293), .C(n7376), .Y(n10077) );
  NAND2X1 U3624 ( .A(arr[1775]), .B(n3294), .Y(n7376) );
  OAI21X1 U3625 ( .A(n5517), .B(n3292), .C(n7377), .Y(n10078) );
  NAND2X1 U3626 ( .A(arr[1776]), .B(n3295), .Y(n7377) );
  OAI21X1 U3627 ( .A(n5519), .B(n3294), .C(n7378), .Y(n10079) );
  NAND2X1 U3628 ( .A(arr[1777]), .B(n3295), .Y(n7378) );
  OAI21X1 U3629 ( .A(n5521), .B(n3294), .C(n7379), .Y(n10080) );
  NAND2X1 U3630 ( .A(arr[1778]), .B(n3295), .Y(n7379) );
  OAI21X1 U3631 ( .A(n5523), .B(n3293), .C(n7380), .Y(n10081) );
  NAND2X1 U3632 ( .A(arr[1779]), .B(n3295), .Y(n7380) );
  OAI21X1 U3633 ( .A(n5525), .B(n3293), .C(n7381), .Y(n10082) );
  NAND2X1 U3634 ( .A(arr[1780]), .B(n3295), .Y(n7381) );
  OAI21X1 U3635 ( .A(n5527), .B(n3293), .C(n7382), .Y(n10083) );
  NAND2X1 U3636 ( .A(arr[1781]), .B(n3295), .Y(n7382) );
  OAI21X1 U3637 ( .A(n5529), .B(n3293), .C(n7383), .Y(n10084) );
  NAND2X1 U3638 ( .A(arr[1782]), .B(n3295), .Y(n7383) );
  OAI21X1 U3639 ( .A(n5531), .B(n3293), .C(n7384), .Y(n10085) );
  NAND2X1 U3640 ( .A(arr[1783]), .B(n3295), .Y(n7384) );
  OAI21X1 U3641 ( .A(n5533), .B(n3293), .C(n7385), .Y(n10086) );
  NAND2X1 U3642 ( .A(arr[1784]), .B(n3295), .Y(n7385) );
  OAI21X1 U3643 ( .A(n5535), .B(n3293), .C(n7386), .Y(n10087) );
  NAND2X1 U3644 ( .A(arr[1785]), .B(n3295), .Y(n7386) );
  OAI21X1 U3645 ( .A(n5537), .B(n3293), .C(n7387), .Y(n10088) );
  NAND2X1 U3646 ( .A(arr[1786]), .B(n3295), .Y(n7387) );
  OAI21X1 U3647 ( .A(n5539), .B(n3293), .C(n7388), .Y(n10089) );
  NAND2X1 U3648 ( .A(arr[1787]), .B(n3295), .Y(n7388) );
  OAI21X1 U3649 ( .A(n5541), .B(n3293), .C(n7389), .Y(n10090) );
  NAND2X1 U3650 ( .A(arr[1788]), .B(n3295), .Y(n7389) );
  OAI21X1 U3651 ( .A(n5543), .B(n3292), .C(n7390), .Y(n10091) );
  NAND2X1 U3652 ( .A(arr[1789]), .B(n3295), .Y(n7390) );
  OAI21X1 U3653 ( .A(n5545), .B(n3292), .C(n7391), .Y(n10092) );
  NAND2X1 U3654 ( .A(arr[1790]), .B(n3295), .Y(n7391) );
  OAI21X1 U3655 ( .A(n5547), .B(n3292), .C(n7392), .Y(n10093) );
  NAND2X1 U3656 ( .A(arr[1791]), .B(n3295), .Y(n7392) );
  OAI21X1 U3657 ( .A(n5549), .B(n3292), .C(n7393), .Y(n10094) );
  NAND2X1 U3658 ( .A(arr[1792]), .B(n3295), .Y(n7393) );
  OAI21X1 U3659 ( .A(n5551), .B(n3292), .C(n7394), .Y(n10095) );
  NAND2X1 U3660 ( .A(arr[1793]), .B(n3296), .Y(n7394) );
  OAI21X1 U3661 ( .A(n5553), .B(n3292), .C(n7395), .Y(n10096) );
  NAND2X1 U3662 ( .A(arr[1794]), .B(n3296), .Y(n7395) );
  OAI21X1 U3663 ( .A(n5555), .B(n3292), .C(n7396), .Y(n10097) );
  NAND2X1 U3664 ( .A(arr[1795]), .B(n3296), .Y(n7396) );
  OAI21X1 U3665 ( .A(n5557), .B(n3292), .C(n7397), .Y(n10098) );
  NAND2X1 U3666 ( .A(arr[1796]), .B(n3296), .Y(n7397) );
  OAI21X1 U3667 ( .A(n5559), .B(n3291), .C(n7398), .Y(n10099) );
  NAND2X1 U3668 ( .A(arr[1797]), .B(n3296), .Y(n7398) );
  OAI21X1 U3669 ( .A(n5561), .B(n3291), .C(n7399), .Y(n10100) );
  NAND2X1 U3670 ( .A(arr[1798]), .B(n3296), .Y(n7399) );
  OAI21X1 U3671 ( .A(n5563), .B(n3291), .C(n7400), .Y(n10101) );
  NAND2X1 U3672 ( .A(arr[1799]), .B(n3296), .Y(n7400) );
  OAI21X1 U3673 ( .A(n5565), .B(n3291), .C(n7401), .Y(n10102) );
  NAND2X1 U3674 ( .A(arr[1800]), .B(n3296), .Y(n7401) );
  OAI21X1 U3675 ( .A(n5567), .B(n3291), .C(n7402), .Y(n10103) );
  NAND2X1 U3676 ( .A(arr[1801]), .B(n3296), .Y(n7402) );
  OAI21X1 U3677 ( .A(n5569), .B(n3291), .C(n7403), .Y(n10104) );
  NAND2X1 U3678 ( .A(arr[1802]), .B(n3294), .Y(n7403) );
  OAI21X1 U3679 ( .A(n5571), .B(n3291), .C(n7404), .Y(n10105) );
  NAND2X1 U3680 ( .A(arr[1803]), .B(n3294), .Y(n7404) );
  NAND2X1 U3681 ( .A(n7278), .B(n5703), .Y(n7363) );
  OAI21X1 U3683 ( .A(n5491), .B(n3285), .C(n7406), .Y(n10106) );
  NAND2X1 U3684 ( .A(arr[1804]), .B(n3288), .Y(n7406) );
  OAI21X1 U3685 ( .A(n5493), .B(n3285), .C(n7407), .Y(n10107) );
  NAND2X1 U3686 ( .A(arr[1805]), .B(n3288), .Y(n7407) );
  OAI21X1 U3687 ( .A(n5495), .B(n3285), .C(n7408), .Y(n10108) );
  NAND2X1 U3688 ( .A(arr[1806]), .B(n3288), .Y(n7408) );
  OAI21X1 U3689 ( .A(n5497), .B(n3285), .C(n7409), .Y(n10109) );
  NAND2X1 U3690 ( .A(arr[1807]), .B(n3288), .Y(n7409) );
  OAI21X1 U3691 ( .A(n5499), .B(n3285), .C(n7410), .Y(n10110) );
  NAND2X1 U3692 ( .A(arr[1808]), .B(n3288), .Y(n7410) );
  OAI21X1 U3693 ( .A(n5501), .B(n3286), .C(n7411), .Y(n10111) );
  NAND2X1 U3694 ( .A(arr[1809]), .B(n3288), .Y(n7411) );
  OAI21X1 U3695 ( .A(n5503), .B(n3286), .C(n7412), .Y(n10112) );
  NAND2X1 U3696 ( .A(arr[1810]), .B(n3288), .Y(n7412) );
  OAI21X1 U3697 ( .A(n5505), .B(n3286), .C(n7413), .Y(n10113) );
  NAND2X1 U3698 ( .A(arr[1811]), .B(n3288), .Y(n7413) );
  OAI21X1 U3699 ( .A(n5507), .B(n3285), .C(n7414), .Y(n10114) );
  NAND2X1 U3700 ( .A(arr[1812]), .B(n3288), .Y(n7414) );
  OAI21X1 U3701 ( .A(n5509), .B(n3286), .C(n7415), .Y(n10115) );
  NAND2X1 U3702 ( .A(arr[1813]), .B(n3288), .Y(n7415) );
  OAI21X1 U3703 ( .A(n5511), .B(n3287), .C(n7416), .Y(n10116) );
  NAND2X1 U3704 ( .A(arr[1814]), .B(n3288), .Y(n7416) );
  OAI21X1 U3705 ( .A(n5513), .B(n3287), .C(n7417), .Y(n10117) );
  NAND2X1 U3706 ( .A(arr[1815]), .B(n3288), .Y(n7417) );
  OAI21X1 U3707 ( .A(n5515), .B(n3287), .C(n7418), .Y(n10118) );
  NAND2X1 U3708 ( .A(arr[1816]), .B(n3288), .Y(n7418) );
  OAI21X1 U3709 ( .A(n5517), .B(n3286), .C(n7419), .Y(n10119) );
  NAND2X1 U3710 ( .A(arr[1817]), .B(n3289), .Y(n7419) );
  OAI21X1 U3711 ( .A(n5519), .B(n3288), .C(n7420), .Y(n10120) );
  NAND2X1 U3712 ( .A(arr[1818]), .B(n3289), .Y(n7420) );
  OAI21X1 U3713 ( .A(n5521), .B(n3288), .C(n7421), .Y(n10121) );
  NAND2X1 U3714 ( .A(arr[1819]), .B(n3289), .Y(n7421) );
  OAI21X1 U3715 ( .A(n5523), .B(n3287), .C(n7422), .Y(n10122) );
  NAND2X1 U3716 ( .A(arr[1820]), .B(n3289), .Y(n7422) );
  OAI21X1 U3717 ( .A(n5525), .B(n3287), .C(n7423), .Y(n10123) );
  NAND2X1 U3718 ( .A(arr[1821]), .B(n3289), .Y(n7423) );
  OAI21X1 U3719 ( .A(n5527), .B(n3287), .C(n7424), .Y(n10124) );
  NAND2X1 U3720 ( .A(arr[1822]), .B(n3289), .Y(n7424) );
  OAI21X1 U3721 ( .A(n5529), .B(n3287), .C(n7425), .Y(n10125) );
  NAND2X1 U3722 ( .A(arr[1823]), .B(n3289), .Y(n7425) );
  OAI21X1 U3723 ( .A(n5531), .B(n3287), .C(n7426), .Y(n10126) );
  NAND2X1 U3724 ( .A(arr[1824]), .B(n3289), .Y(n7426) );
  OAI21X1 U3725 ( .A(n5533), .B(n3287), .C(n7427), .Y(n10127) );
  NAND2X1 U3726 ( .A(arr[1825]), .B(n3289), .Y(n7427) );
  OAI21X1 U3727 ( .A(n5535), .B(n3287), .C(n7428), .Y(n10128) );
  NAND2X1 U3728 ( .A(arr[1826]), .B(n3289), .Y(n7428) );
  OAI21X1 U3729 ( .A(n5537), .B(n3287), .C(n7429), .Y(n10129) );
  NAND2X1 U3730 ( .A(arr[1827]), .B(n3289), .Y(n7429) );
  OAI21X1 U3731 ( .A(n5539), .B(n3287), .C(n7430), .Y(n10130) );
  NAND2X1 U3732 ( .A(arr[1828]), .B(n3289), .Y(n7430) );
  OAI21X1 U3733 ( .A(n5541), .B(n3287), .C(n7431), .Y(n10131) );
  NAND2X1 U3734 ( .A(arr[1829]), .B(n3289), .Y(n7431) );
  OAI21X1 U3735 ( .A(n5543), .B(n3286), .C(n7432), .Y(n10132) );
  NAND2X1 U3736 ( .A(arr[1830]), .B(n3289), .Y(n7432) );
  OAI21X1 U3737 ( .A(n5545), .B(n3286), .C(n7433), .Y(n10133) );
  NAND2X1 U3738 ( .A(arr[1831]), .B(n3289), .Y(n7433) );
  OAI21X1 U3739 ( .A(n5547), .B(n3286), .C(n7434), .Y(n10134) );
  NAND2X1 U3740 ( .A(arr[1832]), .B(n3289), .Y(n7434) );
  OAI21X1 U3741 ( .A(n5549), .B(n3286), .C(n7435), .Y(n10135) );
  NAND2X1 U3742 ( .A(arr[1833]), .B(n3289), .Y(n7435) );
  OAI21X1 U3743 ( .A(n5551), .B(n3286), .C(n7436), .Y(n10136) );
  NAND2X1 U3744 ( .A(arr[1834]), .B(n3290), .Y(n7436) );
  OAI21X1 U3745 ( .A(n5553), .B(n3286), .C(n7437), .Y(n10137) );
  NAND2X1 U3746 ( .A(arr[1835]), .B(n3290), .Y(n7437) );
  OAI21X1 U3747 ( .A(n5555), .B(n3286), .C(n7438), .Y(n10138) );
  NAND2X1 U3748 ( .A(arr[1836]), .B(n3290), .Y(n7438) );
  OAI21X1 U3749 ( .A(n5557), .B(n3286), .C(n7439), .Y(n10139) );
  NAND2X1 U3750 ( .A(arr[1837]), .B(n3290), .Y(n7439) );
  OAI21X1 U3751 ( .A(n5559), .B(n3285), .C(n7440), .Y(n10140) );
  NAND2X1 U3752 ( .A(arr[1838]), .B(n3290), .Y(n7440) );
  OAI21X1 U3753 ( .A(n5561), .B(n3285), .C(n7441), .Y(n10141) );
  NAND2X1 U3754 ( .A(arr[1839]), .B(n3290), .Y(n7441) );
  OAI21X1 U3755 ( .A(n5563), .B(n3285), .C(n7442), .Y(n10142) );
  NAND2X1 U3756 ( .A(arr[1840]), .B(n3290), .Y(n7442) );
  OAI21X1 U3757 ( .A(n5565), .B(n3285), .C(n7443), .Y(n10143) );
  NAND2X1 U3758 ( .A(arr[1841]), .B(n3290), .Y(n7443) );
  OAI21X1 U3759 ( .A(n5567), .B(n3285), .C(n7444), .Y(n10144) );
  NAND2X1 U3760 ( .A(arr[1842]), .B(n3290), .Y(n7444) );
  OAI21X1 U3761 ( .A(n5569), .B(n3285), .C(n7445), .Y(n10145) );
  NAND2X1 U3762 ( .A(arr[1843]), .B(n3288), .Y(n7445) );
  OAI21X1 U3763 ( .A(n5571), .B(n3285), .C(n7446), .Y(n10146) );
  NAND2X1 U3764 ( .A(arr[1844]), .B(n3288), .Y(n7446) );
  NAND2X1 U3765 ( .A(n7447), .B(n5573), .Y(n7405) );
  OAI21X1 U3766 ( .A(n5491), .B(n3279), .C(n7449), .Y(n10147) );
  NAND2X1 U3767 ( .A(arr[1845]), .B(n3282), .Y(n7449) );
  OAI21X1 U3768 ( .A(n5493), .B(n3279), .C(n7450), .Y(n10148) );
  NAND2X1 U3769 ( .A(arr[1846]), .B(n3282), .Y(n7450) );
  OAI21X1 U3770 ( .A(n5495), .B(n3279), .C(n7451), .Y(n10149) );
  NAND2X1 U3771 ( .A(arr[1847]), .B(n3282), .Y(n7451) );
  OAI21X1 U3772 ( .A(n5497), .B(n3279), .C(n7452), .Y(n10150) );
  NAND2X1 U3773 ( .A(arr[1848]), .B(n3282), .Y(n7452) );
  OAI21X1 U3774 ( .A(n5499), .B(n3279), .C(n7453), .Y(n10151) );
  NAND2X1 U3775 ( .A(arr[1849]), .B(n3282), .Y(n7453) );
  OAI21X1 U3776 ( .A(n5501), .B(n3280), .C(n7454), .Y(n10152) );
  NAND2X1 U3777 ( .A(arr[1850]), .B(n3282), .Y(n7454) );
  OAI21X1 U3778 ( .A(n5503), .B(n3280), .C(n7455), .Y(n10153) );
  NAND2X1 U3779 ( .A(arr[1851]), .B(n3282), .Y(n7455) );
  OAI21X1 U3780 ( .A(n5505), .B(n3280), .C(n7456), .Y(n10154) );
  NAND2X1 U3781 ( .A(arr[1852]), .B(n3282), .Y(n7456) );
  OAI21X1 U3782 ( .A(n5507), .B(n3279), .C(n7457), .Y(n10155) );
  NAND2X1 U3783 ( .A(arr[1853]), .B(n3282), .Y(n7457) );
  OAI21X1 U3784 ( .A(n5509), .B(n3280), .C(n7458), .Y(n10156) );
  NAND2X1 U3785 ( .A(arr[1854]), .B(n3282), .Y(n7458) );
  OAI21X1 U3786 ( .A(n5511), .B(n3281), .C(n7459), .Y(n10157) );
  NAND2X1 U3787 ( .A(arr[1855]), .B(n3282), .Y(n7459) );
  OAI21X1 U3788 ( .A(n5513), .B(n3281), .C(n7460), .Y(n10158) );
  NAND2X1 U3789 ( .A(arr[1856]), .B(n3282), .Y(n7460) );
  OAI21X1 U3790 ( .A(n5515), .B(n3281), .C(n7461), .Y(n10159) );
  NAND2X1 U3791 ( .A(arr[1857]), .B(n3282), .Y(n7461) );
  OAI21X1 U3792 ( .A(n5517), .B(n3280), .C(n7462), .Y(n10160) );
  NAND2X1 U3793 ( .A(arr[1858]), .B(n3283), .Y(n7462) );
  OAI21X1 U3794 ( .A(n5519), .B(n3282), .C(n7463), .Y(n10161) );
  NAND2X1 U3795 ( .A(arr[1859]), .B(n3283), .Y(n7463) );
  OAI21X1 U3796 ( .A(n5521), .B(n3282), .C(n7464), .Y(n10162) );
  NAND2X1 U3797 ( .A(arr[1860]), .B(n3283), .Y(n7464) );
  OAI21X1 U3798 ( .A(n5523), .B(n3281), .C(n7465), .Y(n10163) );
  NAND2X1 U3799 ( .A(arr[1861]), .B(n3283), .Y(n7465) );
  OAI21X1 U3800 ( .A(n5525), .B(n3281), .C(n7466), .Y(n10164) );
  NAND2X1 U3801 ( .A(arr[1862]), .B(n3283), .Y(n7466) );
  OAI21X1 U3802 ( .A(n5527), .B(n3281), .C(n7467), .Y(n10165) );
  NAND2X1 U3803 ( .A(arr[1863]), .B(n3283), .Y(n7467) );
  OAI21X1 U3804 ( .A(n5529), .B(n3281), .C(n7468), .Y(n10166) );
  NAND2X1 U3805 ( .A(arr[1864]), .B(n3283), .Y(n7468) );
  OAI21X1 U3806 ( .A(n5531), .B(n3281), .C(n7469), .Y(n10167) );
  NAND2X1 U3807 ( .A(arr[1865]), .B(n3283), .Y(n7469) );
  OAI21X1 U3808 ( .A(n5533), .B(n3281), .C(n7470), .Y(n10168) );
  NAND2X1 U3809 ( .A(arr[1866]), .B(n3283), .Y(n7470) );
  OAI21X1 U3810 ( .A(n5535), .B(n3281), .C(n7471), .Y(n10169) );
  NAND2X1 U3811 ( .A(arr[1867]), .B(n3283), .Y(n7471) );
  OAI21X1 U3812 ( .A(n5537), .B(n3281), .C(n7472), .Y(n10170) );
  NAND2X1 U3813 ( .A(arr[1868]), .B(n3283), .Y(n7472) );
  OAI21X1 U3814 ( .A(n5539), .B(n3281), .C(n7473), .Y(n10171) );
  NAND2X1 U3815 ( .A(arr[1869]), .B(n3283), .Y(n7473) );
  OAI21X1 U3816 ( .A(n5541), .B(n3281), .C(n7474), .Y(n10172) );
  NAND2X1 U3817 ( .A(arr[1870]), .B(n3283), .Y(n7474) );
  OAI21X1 U3818 ( .A(n5543), .B(n3280), .C(n7475), .Y(n10173) );
  NAND2X1 U3819 ( .A(arr[1871]), .B(n3283), .Y(n7475) );
  OAI21X1 U3820 ( .A(n5545), .B(n3280), .C(n7476), .Y(n10174) );
  NAND2X1 U3821 ( .A(arr[1872]), .B(n3283), .Y(n7476) );
  OAI21X1 U3822 ( .A(n5547), .B(n3280), .C(n7477), .Y(n10175) );
  NAND2X1 U3823 ( .A(arr[1873]), .B(n3283), .Y(n7477) );
  OAI21X1 U3824 ( .A(n5549), .B(n3280), .C(n7478), .Y(n10176) );
  NAND2X1 U3825 ( .A(arr[1874]), .B(n3283), .Y(n7478) );
  OAI21X1 U3826 ( .A(n5551), .B(n3280), .C(n7479), .Y(n10177) );
  NAND2X1 U3827 ( .A(arr[1875]), .B(n3284), .Y(n7479) );
  OAI21X1 U3828 ( .A(n5553), .B(n3280), .C(n7480), .Y(n10178) );
  NAND2X1 U3829 ( .A(arr[1876]), .B(n3284), .Y(n7480) );
  OAI21X1 U3830 ( .A(n5555), .B(n3280), .C(n7481), .Y(n10179) );
  NAND2X1 U3831 ( .A(arr[1877]), .B(n3284), .Y(n7481) );
  OAI21X1 U3832 ( .A(n5557), .B(n3280), .C(n7482), .Y(n10180) );
  NAND2X1 U3833 ( .A(arr[1878]), .B(n3284), .Y(n7482) );
  OAI21X1 U3834 ( .A(n5559), .B(n3279), .C(n7483), .Y(n10181) );
  NAND2X1 U3835 ( .A(arr[1879]), .B(n3284), .Y(n7483) );
  OAI21X1 U3836 ( .A(n5561), .B(n3279), .C(n7484), .Y(n10182) );
  NAND2X1 U3837 ( .A(arr[1880]), .B(n3284), .Y(n7484) );
  OAI21X1 U3838 ( .A(n5563), .B(n3279), .C(n7485), .Y(n10183) );
  NAND2X1 U3839 ( .A(arr[1881]), .B(n3284), .Y(n7485) );
  OAI21X1 U3840 ( .A(n5565), .B(n3279), .C(n7486), .Y(n10184) );
  NAND2X1 U3841 ( .A(arr[1882]), .B(n3284), .Y(n7486) );
  OAI21X1 U3842 ( .A(n5567), .B(n3279), .C(n7487), .Y(n10185) );
  NAND2X1 U3843 ( .A(arr[1883]), .B(n3284), .Y(n7487) );
  OAI21X1 U3844 ( .A(n5569), .B(n3279), .C(n7488), .Y(n10186) );
  NAND2X1 U3845 ( .A(arr[1884]), .B(n3282), .Y(n7488) );
  OAI21X1 U3846 ( .A(n5571), .B(n3279), .C(n7489), .Y(n10187) );
  NAND2X1 U3847 ( .A(arr[1885]), .B(n3282), .Y(n7489) );
  NAND2X1 U3848 ( .A(n7447), .B(n5617), .Y(n7448) );
  OAI21X1 U3849 ( .A(n5491), .B(n3273), .C(n7491), .Y(n10188) );
  NAND2X1 U3850 ( .A(arr[1886]), .B(n3276), .Y(n7491) );
  OAI21X1 U3851 ( .A(n5493), .B(n3273), .C(n7492), .Y(n10189) );
  NAND2X1 U3852 ( .A(arr[1887]), .B(n3276), .Y(n7492) );
  OAI21X1 U3853 ( .A(n5495), .B(n3273), .C(n7493), .Y(n10190) );
  NAND2X1 U3854 ( .A(arr[1888]), .B(n3276), .Y(n7493) );
  OAI21X1 U3855 ( .A(n5497), .B(n3273), .C(n7494), .Y(n10191) );
  NAND2X1 U3856 ( .A(arr[1889]), .B(n3276), .Y(n7494) );
  OAI21X1 U3857 ( .A(n5499), .B(n3273), .C(n7495), .Y(n10192) );
  NAND2X1 U3858 ( .A(arr[1890]), .B(n3276), .Y(n7495) );
  OAI21X1 U3859 ( .A(n5501), .B(n3274), .C(n7496), .Y(n10193) );
  NAND2X1 U3860 ( .A(arr[1891]), .B(n3276), .Y(n7496) );
  OAI21X1 U3861 ( .A(n5503), .B(n3274), .C(n7497), .Y(n10194) );
  NAND2X1 U3862 ( .A(arr[1892]), .B(n3276), .Y(n7497) );
  OAI21X1 U3863 ( .A(n5505), .B(n3274), .C(n7498), .Y(n10195) );
  NAND2X1 U3864 ( .A(arr[1893]), .B(n3276), .Y(n7498) );
  OAI21X1 U3865 ( .A(n5507), .B(n3273), .C(n7499), .Y(n10196) );
  NAND2X1 U3866 ( .A(arr[1894]), .B(n3276), .Y(n7499) );
  OAI21X1 U3867 ( .A(n5509), .B(n3274), .C(n7500), .Y(n10197) );
  NAND2X1 U3868 ( .A(arr[1895]), .B(n3276), .Y(n7500) );
  OAI21X1 U3869 ( .A(n5511), .B(n3275), .C(n7501), .Y(n10198) );
  NAND2X1 U3870 ( .A(arr[1896]), .B(n3276), .Y(n7501) );
  OAI21X1 U3871 ( .A(n5513), .B(n3275), .C(n7502), .Y(n10199) );
  NAND2X1 U3872 ( .A(arr[1897]), .B(n3276), .Y(n7502) );
  OAI21X1 U3873 ( .A(n5515), .B(n3275), .C(n7503), .Y(n10200) );
  NAND2X1 U3874 ( .A(arr[1898]), .B(n3276), .Y(n7503) );
  OAI21X1 U3875 ( .A(n5517), .B(n3274), .C(n7504), .Y(n10201) );
  NAND2X1 U3876 ( .A(arr[1899]), .B(n3277), .Y(n7504) );
  OAI21X1 U3877 ( .A(n5519), .B(n3276), .C(n7505), .Y(n10202) );
  NAND2X1 U3878 ( .A(arr[1900]), .B(n3277), .Y(n7505) );
  OAI21X1 U3879 ( .A(n5521), .B(n3276), .C(n7506), .Y(n10203) );
  NAND2X1 U3880 ( .A(arr[1901]), .B(n3277), .Y(n7506) );
  OAI21X1 U3881 ( .A(n5523), .B(n3275), .C(n7507), .Y(n10204) );
  NAND2X1 U3882 ( .A(arr[1902]), .B(n3277), .Y(n7507) );
  OAI21X1 U3883 ( .A(n5525), .B(n3275), .C(n7508), .Y(n10205) );
  NAND2X1 U3884 ( .A(arr[1903]), .B(n3277), .Y(n7508) );
  OAI21X1 U3885 ( .A(n5527), .B(n3275), .C(n7509), .Y(n10206) );
  NAND2X1 U3886 ( .A(arr[1904]), .B(n3277), .Y(n7509) );
  OAI21X1 U3887 ( .A(n5529), .B(n3275), .C(n7510), .Y(n10207) );
  NAND2X1 U3888 ( .A(arr[1905]), .B(n3277), .Y(n7510) );
  OAI21X1 U3889 ( .A(n5531), .B(n3275), .C(n7511), .Y(n10208) );
  NAND2X1 U3890 ( .A(arr[1906]), .B(n3277), .Y(n7511) );
  OAI21X1 U3891 ( .A(n5533), .B(n3275), .C(n7512), .Y(n10209) );
  NAND2X1 U3892 ( .A(arr[1907]), .B(n3277), .Y(n7512) );
  OAI21X1 U3893 ( .A(n5535), .B(n3275), .C(n7513), .Y(n10210) );
  NAND2X1 U3894 ( .A(arr[1908]), .B(n3277), .Y(n7513) );
  OAI21X1 U3895 ( .A(n5537), .B(n3275), .C(n7514), .Y(n10211) );
  NAND2X1 U3896 ( .A(arr[1909]), .B(n3277), .Y(n7514) );
  OAI21X1 U3897 ( .A(n5539), .B(n3275), .C(n7515), .Y(n10212) );
  NAND2X1 U3898 ( .A(arr[1910]), .B(n3277), .Y(n7515) );
  OAI21X1 U3899 ( .A(n5541), .B(n3275), .C(n7516), .Y(n10213) );
  NAND2X1 U3900 ( .A(arr[1911]), .B(n3277), .Y(n7516) );
  OAI21X1 U3901 ( .A(n5543), .B(n3274), .C(n7517), .Y(n10214) );
  NAND2X1 U3902 ( .A(arr[1912]), .B(n3277), .Y(n7517) );
  OAI21X1 U3903 ( .A(n5545), .B(n3274), .C(n7518), .Y(n10215) );
  NAND2X1 U3904 ( .A(arr[1913]), .B(n3277), .Y(n7518) );
  OAI21X1 U3905 ( .A(n5547), .B(n3274), .C(n7519), .Y(n10216) );
  NAND2X1 U3906 ( .A(arr[1914]), .B(n3277), .Y(n7519) );
  OAI21X1 U3907 ( .A(n5549), .B(n3274), .C(n7520), .Y(n10217) );
  NAND2X1 U3908 ( .A(arr[1915]), .B(n3277), .Y(n7520) );
  OAI21X1 U3909 ( .A(n5551), .B(n3274), .C(n7521), .Y(n10218) );
  NAND2X1 U3910 ( .A(arr[1916]), .B(n3278), .Y(n7521) );
  OAI21X1 U3911 ( .A(n5553), .B(n3274), .C(n7522), .Y(n10219) );
  NAND2X1 U3912 ( .A(arr[1917]), .B(n3278), .Y(n7522) );
  OAI21X1 U3913 ( .A(n5555), .B(n3274), .C(n7523), .Y(n10220) );
  NAND2X1 U3914 ( .A(arr[1918]), .B(n3278), .Y(n7523) );
  OAI21X1 U3915 ( .A(n5557), .B(n3274), .C(n7524), .Y(n10221) );
  NAND2X1 U3916 ( .A(arr[1919]), .B(n3278), .Y(n7524) );
  OAI21X1 U3917 ( .A(n5559), .B(n3273), .C(n7525), .Y(n10222) );
  NAND2X1 U3918 ( .A(arr[1920]), .B(n3278), .Y(n7525) );
  OAI21X1 U3919 ( .A(n5561), .B(n3273), .C(n7526), .Y(n10223) );
  NAND2X1 U3920 ( .A(arr[1921]), .B(n3278), .Y(n7526) );
  OAI21X1 U3921 ( .A(n5563), .B(n3273), .C(n7527), .Y(n10224) );
  NAND2X1 U3922 ( .A(arr[1922]), .B(n3278), .Y(n7527) );
  OAI21X1 U3923 ( .A(n5565), .B(n3273), .C(n7528), .Y(n10225) );
  NAND2X1 U3924 ( .A(arr[1923]), .B(n3278), .Y(n7528) );
  OAI21X1 U3925 ( .A(n5567), .B(n3273), .C(n7529), .Y(n10226) );
  NAND2X1 U3926 ( .A(arr[1924]), .B(n3278), .Y(n7529) );
  OAI21X1 U3927 ( .A(n5569), .B(n3273), .C(n7530), .Y(n10227) );
  NAND2X1 U3928 ( .A(arr[1925]), .B(n3276), .Y(n7530) );
  OAI21X1 U3929 ( .A(n5571), .B(n3273), .C(n7531), .Y(n10228) );
  NAND2X1 U3930 ( .A(arr[1926]), .B(n3276), .Y(n7531) );
  NAND2X1 U3931 ( .A(n7447), .B(n5660), .Y(n7490) );
  OAI21X1 U3932 ( .A(n5491), .B(n3267), .C(n7533), .Y(n10229) );
  NAND2X1 U3933 ( .A(arr[1927]), .B(n3270), .Y(n7533) );
  OAI21X1 U3934 ( .A(n5493), .B(n3267), .C(n7534), .Y(n10230) );
  NAND2X1 U3935 ( .A(arr[1928]), .B(n3270), .Y(n7534) );
  OAI21X1 U3936 ( .A(n5495), .B(n3267), .C(n7535), .Y(n10231) );
  NAND2X1 U3937 ( .A(arr[1929]), .B(n3270), .Y(n7535) );
  OAI21X1 U3938 ( .A(n5497), .B(n3267), .C(n7536), .Y(n10232) );
  NAND2X1 U3939 ( .A(arr[1930]), .B(n3270), .Y(n7536) );
  OAI21X1 U3940 ( .A(n5499), .B(n3267), .C(n7537), .Y(n10233) );
  NAND2X1 U3941 ( .A(arr[1931]), .B(n3270), .Y(n7537) );
  OAI21X1 U3942 ( .A(n5501), .B(n3268), .C(n7538), .Y(n10234) );
  NAND2X1 U3943 ( .A(arr[1932]), .B(n3270), .Y(n7538) );
  OAI21X1 U3944 ( .A(n5503), .B(n3268), .C(n7539), .Y(n10235) );
  NAND2X1 U3945 ( .A(arr[1933]), .B(n3270), .Y(n7539) );
  OAI21X1 U3946 ( .A(n5505), .B(n3268), .C(n7540), .Y(n10236) );
  NAND2X1 U3947 ( .A(arr[1934]), .B(n3270), .Y(n7540) );
  OAI21X1 U3948 ( .A(n5507), .B(n3267), .C(n7541), .Y(n10237) );
  NAND2X1 U3949 ( .A(arr[1935]), .B(n3270), .Y(n7541) );
  OAI21X1 U3950 ( .A(n5509), .B(n3268), .C(n7542), .Y(n10238) );
  NAND2X1 U3951 ( .A(arr[1936]), .B(n3270), .Y(n7542) );
  OAI21X1 U3952 ( .A(n5511), .B(n3269), .C(n7543), .Y(n10239) );
  NAND2X1 U3953 ( .A(arr[1937]), .B(n3270), .Y(n7543) );
  OAI21X1 U3954 ( .A(n5513), .B(n3269), .C(n7544), .Y(n10240) );
  NAND2X1 U3955 ( .A(arr[1938]), .B(n3270), .Y(n7544) );
  OAI21X1 U3956 ( .A(n5515), .B(n3269), .C(n7545), .Y(n10241) );
  NAND2X1 U3957 ( .A(arr[1939]), .B(n3270), .Y(n7545) );
  OAI21X1 U3958 ( .A(n5517), .B(n3268), .C(n7546), .Y(n10242) );
  NAND2X1 U3959 ( .A(arr[1940]), .B(n3271), .Y(n7546) );
  OAI21X1 U3960 ( .A(n5519), .B(n3270), .C(n7547), .Y(n10243) );
  NAND2X1 U3961 ( .A(arr[1941]), .B(n3271), .Y(n7547) );
  OAI21X1 U3962 ( .A(n5521), .B(n3270), .C(n7548), .Y(n10244) );
  NAND2X1 U3963 ( .A(arr[1942]), .B(n3271), .Y(n7548) );
  OAI21X1 U3964 ( .A(n5523), .B(n3269), .C(n7549), .Y(n10245) );
  NAND2X1 U3965 ( .A(arr[1943]), .B(n3271), .Y(n7549) );
  OAI21X1 U3966 ( .A(n5525), .B(n3269), .C(n7550), .Y(n10246) );
  NAND2X1 U3967 ( .A(arr[1944]), .B(n3271), .Y(n7550) );
  OAI21X1 U3968 ( .A(n5527), .B(n3269), .C(n7551), .Y(n10247) );
  NAND2X1 U3969 ( .A(arr[1945]), .B(n3271), .Y(n7551) );
  OAI21X1 U3970 ( .A(n5529), .B(n3269), .C(n7552), .Y(n10248) );
  NAND2X1 U3971 ( .A(arr[1946]), .B(n3271), .Y(n7552) );
  OAI21X1 U3972 ( .A(n5531), .B(n3269), .C(n7553), .Y(n10249) );
  NAND2X1 U3973 ( .A(arr[1947]), .B(n3271), .Y(n7553) );
  OAI21X1 U3974 ( .A(n5533), .B(n3269), .C(n7554), .Y(n10250) );
  NAND2X1 U3975 ( .A(arr[1948]), .B(n3271), .Y(n7554) );
  OAI21X1 U3976 ( .A(n5535), .B(n3269), .C(n7555), .Y(n10251) );
  NAND2X1 U3977 ( .A(arr[1949]), .B(n3271), .Y(n7555) );
  OAI21X1 U3978 ( .A(n5537), .B(n3269), .C(n7556), .Y(n10252) );
  NAND2X1 U3979 ( .A(arr[1950]), .B(n3271), .Y(n7556) );
  OAI21X1 U3980 ( .A(n5539), .B(n3269), .C(n7557), .Y(n10253) );
  NAND2X1 U3981 ( .A(arr[1951]), .B(n3271), .Y(n7557) );
  OAI21X1 U3982 ( .A(n5541), .B(n3269), .C(n7558), .Y(n10254) );
  NAND2X1 U3983 ( .A(arr[1952]), .B(n3271), .Y(n7558) );
  OAI21X1 U3984 ( .A(n5543), .B(n3268), .C(n7559), .Y(n10255) );
  NAND2X1 U3985 ( .A(arr[1953]), .B(n3271), .Y(n7559) );
  OAI21X1 U3986 ( .A(n5545), .B(n3268), .C(n7560), .Y(n10256) );
  NAND2X1 U3987 ( .A(arr[1954]), .B(n3271), .Y(n7560) );
  OAI21X1 U3988 ( .A(n5547), .B(n3268), .C(n7561), .Y(n10257) );
  NAND2X1 U3989 ( .A(arr[1955]), .B(n3271), .Y(n7561) );
  OAI21X1 U3990 ( .A(n5549), .B(n3268), .C(n7562), .Y(n10258) );
  NAND2X1 U3991 ( .A(arr[1956]), .B(n3271), .Y(n7562) );
  OAI21X1 U3992 ( .A(n5551), .B(n3268), .C(n7563), .Y(n10259) );
  NAND2X1 U3993 ( .A(arr[1957]), .B(n3272), .Y(n7563) );
  OAI21X1 U3994 ( .A(n5553), .B(n3268), .C(n7564), .Y(n10260) );
  NAND2X1 U3995 ( .A(arr[1958]), .B(n3272), .Y(n7564) );
  OAI21X1 U3996 ( .A(n5555), .B(n3268), .C(n7565), .Y(n10261) );
  NAND2X1 U3997 ( .A(arr[1959]), .B(n3272), .Y(n7565) );
  OAI21X1 U3998 ( .A(n5557), .B(n3268), .C(n7566), .Y(n10262) );
  NAND2X1 U3999 ( .A(arr[1960]), .B(n3272), .Y(n7566) );
  OAI21X1 U4000 ( .A(n5559), .B(n3267), .C(n7567), .Y(n10263) );
  NAND2X1 U4001 ( .A(arr[1961]), .B(n3272), .Y(n7567) );
  OAI21X1 U4002 ( .A(n5561), .B(n3267), .C(n7568), .Y(n10264) );
  NAND2X1 U4003 ( .A(arr[1962]), .B(n3272), .Y(n7568) );
  OAI21X1 U4004 ( .A(n5563), .B(n3267), .C(n7569), .Y(n10265) );
  NAND2X1 U4005 ( .A(arr[1963]), .B(n3272), .Y(n7569) );
  OAI21X1 U4006 ( .A(n5565), .B(n3267), .C(n7570), .Y(n10266) );
  NAND2X1 U4007 ( .A(arr[1964]), .B(n3272), .Y(n7570) );
  OAI21X1 U4008 ( .A(n5567), .B(n3267), .C(n7571), .Y(n10267) );
  NAND2X1 U4009 ( .A(arr[1965]), .B(n3272), .Y(n7571) );
  OAI21X1 U4010 ( .A(n5569), .B(n3267), .C(n7572), .Y(n10268) );
  NAND2X1 U4011 ( .A(arr[1966]), .B(n3270), .Y(n7572) );
  OAI21X1 U4012 ( .A(n5571), .B(n3267), .C(n7573), .Y(n10269) );
  NAND2X1 U4013 ( .A(arr[1967]), .B(n3270), .Y(n7573) );
  NAND2X1 U4014 ( .A(n7447), .B(n5703), .Y(n7532) );
  AND2X1 U4016 ( .A(n7574), .B(n6217), .Y(n7066) );
  OAI21X1 U4017 ( .A(n5491), .B(n3261), .C(n7576), .Y(n10270) );
  NAND2X1 U4018 ( .A(arr[1968]), .B(n3264), .Y(n7576) );
  OAI21X1 U4019 ( .A(n5493), .B(n3261), .C(n7577), .Y(n10271) );
  NAND2X1 U4020 ( .A(arr[1969]), .B(n3264), .Y(n7577) );
  OAI21X1 U4021 ( .A(n5495), .B(n3261), .C(n7578), .Y(n10272) );
  NAND2X1 U4022 ( .A(arr[1970]), .B(n3264), .Y(n7578) );
  OAI21X1 U4023 ( .A(n5497), .B(n3261), .C(n7579), .Y(n10273) );
  NAND2X1 U4024 ( .A(arr[1971]), .B(n3264), .Y(n7579) );
  OAI21X1 U4025 ( .A(n5499), .B(n3261), .C(n7580), .Y(n10274) );
  NAND2X1 U4026 ( .A(arr[1972]), .B(n3264), .Y(n7580) );
  OAI21X1 U4027 ( .A(n5501), .B(n3262), .C(n7581), .Y(n10275) );
  NAND2X1 U4028 ( .A(arr[1973]), .B(n3264), .Y(n7581) );
  OAI21X1 U4029 ( .A(n5503), .B(n3262), .C(n7582), .Y(n10276) );
  NAND2X1 U4030 ( .A(arr[1974]), .B(n3264), .Y(n7582) );
  OAI21X1 U4031 ( .A(n5505), .B(n3262), .C(n7583), .Y(n10277) );
  NAND2X1 U4032 ( .A(arr[1975]), .B(n3264), .Y(n7583) );
  OAI21X1 U4033 ( .A(n5507), .B(n3261), .C(n7584), .Y(n10278) );
  NAND2X1 U4034 ( .A(arr[1976]), .B(n3264), .Y(n7584) );
  OAI21X1 U4035 ( .A(n5509), .B(n3262), .C(n7585), .Y(n10279) );
  NAND2X1 U4036 ( .A(arr[1977]), .B(n3264), .Y(n7585) );
  OAI21X1 U4037 ( .A(n5511), .B(n3263), .C(n7586), .Y(n10280) );
  NAND2X1 U4038 ( .A(arr[1978]), .B(n3264), .Y(n7586) );
  OAI21X1 U4039 ( .A(n5513), .B(n3263), .C(n7587), .Y(n10281) );
  NAND2X1 U4040 ( .A(arr[1979]), .B(n3264), .Y(n7587) );
  OAI21X1 U4041 ( .A(n5515), .B(n3263), .C(n7588), .Y(n10282) );
  NAND2X1 U4042 ( .A(arr[1980]), .B(n3264), .Y(n7588) );
  OAI21X1 U4043 ( .A(n5517), .B(n3262), .C(n7589), .Y(n10283) );
  NAND2X1 U4044 ( .A(arr[1981]), .B(n3265), .Y(n7589) );
  OAI21X1 U4045 ( .A(n5519), .B(n3264), .C(n7590), .Y(n10284) );
  NAND2X1 U4046 ( .A(arr[1982]), .B(n3265), .Y(n7590) );
  OAI21X1 U4047 ( .A(n5521), .B(n3264), .C(n7591), .Y(n10285) );
  NAND2X1 U4048 ( .A(arr[1983]), .B(n3265), .Y(n7591) );
  OAI21X1 U4049 ( .A(n5523), .B(n3263), .C(n7592), .Y(n10286) );
  NAND2X1 U4050 ( .A(arr[1984]), .B(n3265), .Y(n7592) );
  OAI21X1 U4051 ( .A(n5525), .B(n3263), .C(n7593), .Y(n10287) );
  NAND2X1 U4052 ( .A(arr[1985]), .B(n3265), .Y(n7593) );
  OAI21X1 U4053 ( .A(n5527), .B(n3263), .C(n7594), .Y(n10288) );
  NAND2X1 U4054 ( .A(arr[1986]), .B(n3265), .Y(n7594) );
  OAI21X1 U4055 ( .A(n5529), .B(n3263), .C(n7595), .Y(n10289) );
  NAND2X1 U4056 ( .A(arr[1987]), .B(n3265), .Y(n7595) );
  OAI21X1 U4057 ( .A(n5531), .B(n3263), .C(n7596), .Y(n10290) );
  NAND2X1 U4058 ( .A(arr[1988]), .B(n3265), .Y(n7596) );
  OAI21X1 U4059 ( .A(n5533), .B(n3263), .C(n7597), .Y(n10291) );
  NAND2X1 U4060 ( .A(arr[1989]), .B(n3265), .Y(n7597) );
  OAI21X1 U4061 ( .A(n5535), .B(n3263), .C(n7598), .Y(n10292) );
  NAND2X1 U4062 ( .A(arr[1990]), .B(n3265), .Y(n7598) );
  OAI21X1 U4063 ( .A(n5537), .B(n3263), .C(n7599), .Y(n10293) );
  NAND2X1 U4064 ( .A(arr[1991]), .B(n3265), .Y(n7599) );
  OAI21X1 U4065 ( .A(n5539), .B(n3263), .C(n7600), .Y(n10294) );
  NAND2X1 U4066 ( .A(arr[1992]), .B(n3265), .Y(n7600) );
  OAI21X1 U4067 ( .A(n5541), .B(n3263), .C(n7601), .Y(n10295) );
  NAND2X1 U4068 ( .A(arr[1993]), .B(n3265), .Y(n7601) );
  OAI21X1 U4069 ( .A(n5543), .B(n3262), .C(n7602), .Y(n10296) );
  NAND2X1 U4070 ( .A(arr[1994]), .B(n3265), .Y(n7602) );
  OAI21X1 U4071 ( .A(n5545), .B(n3262), .C(n7603), .Y(n10297) );
  NAND2X1 U4072 ( .A(arr[1995]), .B(n3265), .Y(n7603) );
  OAI21X1 U4073 ( .A(n5547), .B(n3262), .C(n7604), .Y(n10298) );
  NAND2X1 U4074 ( .A(arr[1996]), .B(n3265), .Y(n7604) );
  OAI21X1 U4075 ( .A(n5549), .B(n3262), .C(n7605), .Y(n10299) );
  NAND2X1 U4076 ( .A(arr[1997]), .B(n3265), .Y(n7605) );
  OAI21X1 U4077 ( .A(n5551), .B(n3262), .C(n7606), .Y(n10300) );
  NAND2X1 U4078 ( .A(arr[1998]), .B(n3266), .Y(n7606) );
  OAI21X1 U4079 ( .A(n5553), .B(n3262), .C(n7607), .Y(n10301) );
  NAND2X1 U4080 ( .A(arr[1999]), .B(n3266), .Y(n7607) );
  OAI21X1 U4081 ( .A(n5555), .B(n3262), .C(n7608), .Y(n10302) );
  NAND2X1 U4082 ( .A(arr[2000]), .B(n3266), .Y(n7608) );
  OAI21X1 U4083 ( .A(n5557), .B(n3262), .C(n7609), .Y(n10303) );
  NAND2X1 U4084 ( .A(arr[2001]), .B(n3266), .Y(n7609) );
  OAI21X1 U4085 ( .A(n5559), .B(n3261), .C(n7610), .Y(n10304) );
  NAND2X1 U4086 ( .A(arr[2002]), .B(n3266), .Y(n7610) );
  OAI21X1 U4087 ( .A(n5561), .B(n3261), .C(n7611), .Y(n10305) );
  NAND2X1 U4088 ( .A(arr[2003]), .B(n3266), .Y(n7611) );
  OAI21X1 U4089 ( .A(n5563), .B(n3261), .C(n7612), .Y(n10306) );
  NAND2X1 U4090 ( .A(arr[2004]), .B(n3266), .Y(n7612) );
  OAI21X1 U4091 ( .A(n5565), .B(n3261), .C(n7613), .Y(n10307) );
  NAND2X1 U4092 ( .A(arr[2005]), .B(n3266), .Y(n7613) );
  OAI21X1 U4093 ( .A(n5567), .B(n3261), .C(n7614), .Y(n10308) );
  NAND2X1 U4094 ( .A(arr[2006]), .B(n3266), .Y(n7614) );
  OAI21X1 U4095 ( .A(n5569), .B(n3261), .C(n7615), .Y(n10309) );
  NAND2X1 U4096 ( .A(arr[2007]), .B(n3264), .Y(n7615) );
  OAI21X1 U4097 ( .A(n5571), .B(n3261), .C(n7616), .Y(n10310) );
  NAND2X1 U4098 ( .A(arr[2008]), .B(n3264), .Y(n7616) );
  NAND2X1 U4099 ( .A(n7617), .B(n5573), .Y(n7575) );
  OAI21X1 U4100 ( .A(n5491), .B(n3255), .C(n7619), .Y(n10311) );
  NAND2X1 U4101 ( .A(arr[2009]), .B(n3258), .Y(n7619) );
  OAI21X1 U4102 ( .A(n5493), .B(n3255), .C(n7620), .Y(n10312) );
  NAND2X1 U4103 ( .A(arr[2010]), .B(n3258), .Y(n7620) );
  OAI21X1 U4104 ( .A(n5495), .B(n3255), .C(n7621), .Y(n10313) );
  NAND2X1 U4105 ( .A(arr[2011]), .B(n3258), .Y(n7621) );
  OAI21X1 U4106 ( .A(n5497), .B(n3255), .C(n7622), .Y(n10314) );
  NAND2X1 U4107 ( .A(arr[2012]), .B(n3258), .Y(n7622) );
  OAI21X1 U4108 ( .A(n5499), .B(n3255), .C(n7623), .Y(n10315) );
  NAND2X1 U4109 ( .A(arr[2013]), .B(n3258), .Y(n7623) );
  OAI21X1 U4110 ( .A(n5501), .B(n3256), .C(n7624), .Y(n10316) );
  NAND2X1 U4111 ( .A(arr[2014]), .B(n3258), .Y(n7624) );
  OAI21X1 U4112 ( .A(n5503), .B(n3256), .C(n7625), .Y(n10317) );
  NAND2X1 U4113 ( .A(arr[2015]), .B(n3258), .Y(n7625) );
  OAI21X1 U4114 ( .A(n5505), .B(n3256), .C(n7626), .Y(n10318) );
  NAND2X1 U4115 ( .A(arr[2016]), .B(n3258), .Y(n7626) );
  OAI21X1 U4116 ( .A(n5507), .B(n3255), .C(n7627), .Y(n10319) );
  NAND2X1 U4117 ( .A(arr[2017]), .B(n3258), .Y(n7627) );
  OAI21X1 U4118 ( .A(n5509), .B(n3256), .C(n7628), .Y(n10320) );
  NAND2X1 U4119 ( .A(arr[2018]), .B(n3258), .Y(n7628) );
  OAI21X1 U4120 ( .A(n5511), .B(n3257), .C(n7629), .Y(n10321) );
  NAND2X1 U4121 ( .A(arr[2019]), .B(n3258), .Y(n7629) );
  OAI21X1 U4122 ( .A(n5513), .B(n3257), .C(n7630), .Y(n10322) );
  NAND2X1 U4123 ( .A(arr[2020]), .B(n3258), .Y(n7630) );
  OAI21X1 U4124 ( .A(n5515), .B(n3257), .C(n7631), .Y(n10323) );
  NAND2X1 U4125 ( .A(arr[2021]), .B(n3258), .Y(n7631) );
  OAI21X1 U4126 ( .A(n5517), .B(n3256), .C(n7632), .Y(n10324) );
  NAND2X1 U4127 ( .A(arr[2022]), .B(n3259), .Y(n7632) );
  OAI21X1 U4128 ( .A(n5519), .B(n3258), .C(n7633), .Y(n10325) );
  NAND2X1 U4129 ( .A(arr[2023]), .B(n3259), .Y(n7633) );
  OAI21X1 U4130 ( .A(n5521), .B(n3258), .C(n7634), .Y(n10326) );
  NAND2X1 U4131 ( .A(arr[2024]), .B(n3259), .Y(n7634) );
  OAI21X1 U4132 ( .A(n5523), .B(n3257), .C(n7635), .Y(n10327) );
  NAND2X1 U4133 ( .A(arr[2025]), .B(n3259), .Y(n7635) );
  OAI21X1 U4134 ( .A(n5525), .B(n3257), .C(n7636), .Y(n10328) );
  NAND2X1 U4135 ( .A(arr[2026]), .B(n3259), .Y(n7636) );
  OAI21X1 U4136 ( .A(n5527), .B(n3257), .C(n7637), .Y(n10329) );
  NAND2X1 U4137 ( .A(arr[2027]), .B(n3259), .Y(n7637) );
  OAI21X1 U4138 ( .A(n5529), .B(n3257), .C(n7638), .Y(n10330) );
  NAND2X1 U4139 ( .A(arr[2028]), .B(n3259), .Y(n7638) );
  OAI21X1 U4140 ( .A(n5531), .B(n3257), .C(n7639), .Y(n10331) );
  NAND2X1 U4141 ( .A(arr[2029]), .B(n3259), .Y(n7639) );
  OAI21X1 U4142 ( .A(n5533), .B(n3257), .C(n7640), .Y(n10332) );
  NAND2X1 U4143 ( .A(arr[2030]), .B(n3259), .Y(n7640) );
  OAI21X1 U4144 ( .A(n5535), .B(n3257), .C(n7641), .Y(n10333) );
  NAND2X1 U4145 ( .A(arr[2031]), .B(n3259), .Y(n7641) );
  OAI21X1 U4146 ( .A(n5537), .B(n3257), .C(n7642), .Y(n10334) );
  NAND2X1 U4147 ( .A(arr[2032]), .B(n3259), .Y(n7642) );
  OAI21X1 U4148 ( .A(n5539), .B(n3257), .C(n7643), .Y(n10335) );
  NAND2X1 U4149 ( .A(arr[2033]), .B(n3259), .Y(n7643) );
  OAI21X1 U4150 ( .A(n5541), .B(n3257), .C(n7644), .Y(n10336) );
  NAND2X1 U4151 ( .A(arr[2034]), .B(n3259), .Y(n7644) );
  OAI21X1 U4152 ( .A(n5543), .B(n3256), .C(n7645), .Y(n10337) );
  NAND2X1 U4153 ( .A(arr[2035]), .B(n3259), .Y(n7645) );
  OAI21X1 U4154 ( .A(n5545), .B(n3256), .C(n7646), .Y(n10338) );
  NAND2X1 U4155 ( .A(arr[2036]), .B(n3259), .Y(n7646) );
  OAI21X1 U4156 ( .A(n5547), .B(n3256), .C(n7647), .Y(n10339) );
  NAND2X1 U4157 ( .A(arr[2037]), .B(n3259), .Y(n7647) );
  OAI21X1 U4158 ( .A(n5549), .B(n3256), .C(n7648), .Y(n10340) );
  NAND2X1 U4159 ( .A(arr[2038]), .B(n3259), .Y(n7648) );
  OAI21X1 U4160 ( .A(n5551), .B(n3256), .C(n7649), .Y(n10341) );
  NAND2X1 U4161 ( .A(arr[2039]), .B(n3260), .Y(n7649) );
  OAI21X1 U4162 ( .A(n5553), .B(n3256), .C(n7650), .Y(n10342) );
  NAND2X1 U4163 ( .A(arr[2040]), .B(n3260), .Y(n7650) );
  OAI21X1 U4164 ( .A(n5555), .B(n3256), .C(n7651), .Y(n10343) );
  NAND2X1 U4165 ( .A(arr[2041]), .B(n3260), .Y(n7651) );
  OAI21X1 U4166 ( .A(n5557), .B(n3256), .C(n7652), .Y(n10344) );
  NAND2X1 U4167 ( .A(arr[2042]), .B(n3260), .Y(n7652) );
  OAI21X1 U4168 ( .A(n5559), .B(n3255), .C(n7653), .Y(n10345) );
  NAND2X1 U4169 ( .A(arr[2043]), .B(n3260), .Y(n7653) );
  OAI21X1 U4170 ( .A(n5561), .B(n3255), .C(n7654), .Y(n10346) );
  NAND2X1 U4171 ( .A(arr[2044]), .B(n3260), .Y(n7654) );
  OAI21X1 U4172 ( .A(n5563), .B(n3255), .C(n7655), .Y(n10347) );
  NAND2X1 U4173 ( .A(arr[2045]), .B(n3260), .Y(n7655) );
  OAI21X1 U4174 ( .A(n5565), .B(n3255), .C(n7656), .Y(n10348) );
  NAND2X1 U4175 ( .A(arr[2046]), .B(n3260), .Y(n7656) );
  OAI21X1 U4176 ( .A(n5567), .B(n3255), .C(n7657), .Y(n10349) );
  NAND2X1 U4177 ( .A(arr[2047]), .B(n3260), .Y(n7657) );
  OAI21X1 U4178 ( .A(n5569), .B(n3255), .C(n7658), .Y(n10350) );
  NAND2X1 U4179 ( .A(arr[2048]), .B(n3258), .Y(n7658) );
  OAI21X1 U4180 ( .A(n5571), .B(n3255), .C(n7659), .Y(n10351) );
  NAND2X1 U4181 ( .A(arr[2049]), .B(n3258), .Y(n7659) );
  NAND2X1 U4182 ( .A(n7617), .B(n5617), .Y(n7618) );
  OAI21X1 U4183 ( .A(n5491), .B(n3249), .C(n7661), .Y(n10352) );
  NAND2X1 U4184 ( .A(arr[2050]), .B(n3252), .Y(n7661) );
  OAI21X1 U4185 ( .A(n5493), .B(n3249), .C(n7662), .Y(n10353) );
  NAND2X1 U4186 ( .A(arr[2051]), .B(n3252), .Y(n7662) );
  OAI21X1 U4187 ( .A(n5495), .B(n3249), .C(n7663), .Y(n10354) );
  NAND2X1 U4188 ( .A(arr[2052]), .B(n3252), .Y(n7663) );
  OAI21X1 U4189 ( .A(n5497), .B(n3249), .C(n7664), .Y(n10355) );
  NAND2X1 U4190 ( .A(arr[2053]), .B(n3252), .Y(n7664) );
  OAI21X1 U4191 ( .A(n5499), .B(n3249), .C(n7665), .Y(n10356) );
  NAND2X1 U4192 ( .A(arr[2054]), .B(n3252), .Y(n7665) );
  OAI21X1 U4193 ( .A(n5501), .B(n3250), .C(n7666), .Y(n10357) );
  NAND2X1 U4194 ( .A(arr[2055]), .B(n3252), .Y(n7666) );
  OAI21X1 U4195 ( .A(n5503), .B(n3250), .C(n7667), .Y(n10358) );
  NAND2X1 U4196 ( .A(arr[2056]), .B(n3252), .Y(n7667) );
  OAI21X1 U4197 ( .A(n5505), .B(n3250), .C(n7668), .Y(n10359) );
  NAND2X1 U4198 ( .A(arr[2057]), .B(n3252), .Y(n7668) );
  OAI21X1 U4199 ( .A(n5507), .B(n3249), .C(n7669), .Y(n10360) );
  NAND2X1 U4200 ( .A(arr[2058]), .B(n3252), .Y(n7669) );
  OAI21X1 U4201 ( .A(n5509), .B(n3250), .C(n7670), .Y(n10361) );
  NAND2X1 U4202 ( .A(arr[2059]), .B(n3252), .Y(n7670) );
  OAI21X1 U4203 ( .A(n5511), .B(n3251), .C(n7671), .Y(n10362) );
  NAND2X1 U4204 ( .A(arr[2060]), .B(n3252), .Y(n7671) );
  OAI21X1 U4205 ( .A(n5513), .B(n3251), .C(n7672), .Y(n10363) );
  NAND2X1 U4206 ( .A(arr[2061]), .B(n3252), .Y(n7672) );
  OAI21X1 U4207 ( .A(n5515), .B(n3251), .C(n7673), .Y(n10364) );
  NAND2X1 U4208 ( .A(arr[2062]), .B(n3252), .Y(n7673) );
  OAI21X1 U4209 ( .A(n5517), .B(n3250), .C(n7674), .Y(n10365) );
  NAND2X1 U4210 ( .A(arr[2063]), .B(n3253), .Y(n7674) );
  OAI21X1 U4211 ( .A(n5519), .B(n3252), .C(n7675), .Y(n10366) );
  NAND2X1 U4212 ( .A(arr[2064]), .B(n3253), .Y(n7675) );
  OAI21X1 U4213 ( .A(n5521), .B(n3252), .C(n7676), .Y(n10367) );
  NAND2X1 U4214 ( .A(arr[2065]), .B(n3253), .Y(n7676) );
  OAI21X1 U4215 ( .A(n5523), .B(n3251), .C(n7677), .Y(n10368) );
  NAND2X1 U4216 ( .A(arr[2066]), .B(n3253), .Y(n7677) );
  OAI21X1 U4217 ( .A(n5525), .B(n3251), .C(n7678), .Y(n10369) );
  NAND2X1 U4218 ( .A(arr[2067]), .B(n3253), .Y(n7678) );
  OAI21X1 U4219 ( .A(n5527), .B(n3251), .C(n7679), .Y(n10370) );
  NAND2X1 U4220 ( .A(arr[2068]), .B(n3253), .Y(n7679) );
  OAI21X1 U4221 ( .A(n5529), .B(n3251), .C(n7680), .Y(n10371) );
  NAND2X1 U4222 ( .A(arr[2069]), .B(n3253), .Y(n7680) );
  OAI21X1 U4223 ( .A(n5531), .B(n3251), .C(n7681), .Y(n10372) );
  NAND2X1 U4224 ( .A(arr[2070]), .B(n3253), .Y(n7681) );
  OAI21X1 U4225 ( .A(n5533), .B(n3251), .C(n7682), .Y(n10373) );
  NAND2X1 U4226 ( .A(arr[2071]), .B(n3253), .Y(n7682) );
  OAI21X1 U4227 ( .A(n5535), .B(n3251), .C(n7683), .Y(n10374) );
  NAND2X1 U4228 ( .A(arr[2072]), .B(n3253), .Y(n7683) );
  OAI21X1 U4229 ( .A(n5537), .B(n3251), .C(n7684), .Y(n10375) );
  NAND2X1 U4230 ( .A(arr[2073]), .B(n3253), .Y(n7684) );
  OAI21X1 U4231 ( .A(n5539), .B(n3251), .C(n7685), .Y(n10376) );
  NAND2X1 U4232 ( .A(arr[2074]), .B(n3253), .Y(n7685) );
  OAI21X1 U4233 ( .A(n5541), .B(n3251), .C(n7686), .Y(n10377) );
  NAND2X1 U4234 ( .A(arr[2075]), .B(n3253), .Y(n7686) );
  OAI21X1 U4235 ( .A(n5543), .B(n3250), .C(n7687), .Y(n10378) );
  NAND2X1 U4236 ( .A(arr[2076]), .B(n3253), .Y(n7687) );
  OAI21X1 U4237 ( .A(n5545), .B(n3250), .C(n7688), .Y(n10379) );
  NAND2X1 U4238 ( .A(arr[2077]), .B(n3253), .Y(n7688) );
  OAI21X1 U4239 ( .A(n5547), .B(n3250), .C(n7689), .Y(n10380) );
  NAND2X1 U4240 ( .A(arr[2078]), .B(n3253), .Y(n7689) );
  OAI21X1 U4241 ( .A(n5549), .B(n3250), .C(n7690), .Y(n10381) );
  NAND2X1 U4242 ( .A(arr[2079]), .B(n3253), .Y(n7690) );
  OAI21X1 U4243 ( .A(n5551), .B(n3250), .C(n7691), .Y(n10382) );
  NAND2X1 U4244 ( .A(arr[2080]), .B(n3254), .Y(n7691) );
  OAI21X1 U4245 ( .A(n5553), .B(n3250), .C(n7692), .Y(n10383) );
  NAND2X1 U4246 ( .A(arr[2081]), .B(n3254), .Y(n7692) );
  OAI21X1 U4247 ( .A(n5555), .B(n3250), .C(n7693), .Y(n10384) );
  NAND2X1 U4248 ( .A(arr[2082]), .B(n3254), .Y(n7693) );
  OAI21X1 U4249 ( .A(n5557), .B(n3250), .C(n7694), .Y(n10385) );
  NAND2X1 U4250 ( .A(arr[2083]), .B(n3254), .Y(n7694) );
  OAI21X1 U4251 ( .A(n5559), .B(n3249), .C(n7695), .Y(n10386) );
  NAND2X1 U4252 ( .A(arr[2084]), .B(n3254), .Y(n7695) );
  OAI21X1 U4253 ( .A(n5561), .B(n3249), .C(n7696), .Y(n10387) );
  NAND2X1 U4254 ( .A(arr[2085]), .B(n3254), .Y(n7696) );
  OAI21X1 U4255 ( .A(n5563), .B(n3249), .C(n7697), .Y(n10388) );
  NAND2X1 U4256 ( .A(arr[2086]), .B(n3254), .Y(n7697) );
  OAI21X1 U4257 ( .A(n5565), .B(n3249), .C(n7698), .Y(n10389) );
  NAND2X1 U4258 ( .A(arr[2087]), .B(n3254), .Y(n7698) );
  OAI21X1 U4259 ( .A(n5567), .B(n3249), .C(n7699), .Y(n10390) );
  NAND2X1 U4260 ( .A(arr[2088]), .B(n3254), .Y(n7699) );
  OAI21X1 U4261 ( .A(n5569), .B(n3249), .C(n7700), .Y(n10391) );
  NAND2X1 U4262 ( .A(arr[2089]), .B(n3252), .Y(n7700) );
  OAI21X1 U4263 ( .A(n5571), .B(n3249), .C(n7701), .Y(n10392) );
  NAND2X1 U4264 ( .A(arr[2090]), .B(n3252), .Y(n7701) );
  NAND2X1 U4265 ( .A(n7617), .B(n5660), .Y(n7660) );
  OAI21X1 U4266 ( .A(n5491), .B(n3243), .C(n7703), .Y(n10393) );
  NAND2X1 U4267 ( .A(arr[2091]), .B(n3246), .Y(n7703) );
  OAI21X1 U4268 ( .A(n5493), .B(n3243), .C(n7704), .Y(n10394) );
  NAND2X1 U4269 ( .A(arr[2092]), .B(n3246), .Y(n7704) );
  OAI21X1 U4270 ( .A(n5495), .B(n3243), .C(n7705), .Y(n10395) );
  NAND2X1 U4271 ( .A(arr[2093]), .B(n3246), .Y(n7705) );
  OAI21X1 U4272 ( .A(n5497), .B(n3243), .C(n7706), .Y(n10396) );
  NAND2X1 U4273 ( .A(arr[2094]), .B(n3246), .Y(n7706) );
  OAI21X1 U4274 ( .A(n5499), .B(n3243), .C(n7707), .Y(n10397) );
  NAND2X1 U4275 ( .A(arr[2095]), .B(n3246), .Y(n7707) );
  OAI21X1 U4276 ( .A(n5501), .B(n3244), .C(n7708), .Y(n10398) );
  NAND2X1 U4277 ( .A(arr[2096]), .B(n3246), .Y(n7708) );
  OAI21X1 U4278 ( .A(n5503), .B(n3244), .C(n7709), .Y(n10399) );
  NAND2X1 U4279 ( .A(arr[2097]), .B(n3246), .Y(n7709) );
  OAI21X1 U4280 ( .A(n5505), .B(n3244), .C(n7710), .Y(n10400) );
  NAND2X1 U4281 ( .A(arr[2098]), .B(n3246), .Y(n7710) );
  OAI21X1 U4282 ( .A(n5507), .B(n3243), .C(n7711), .Y(n10401) );
  NAND2X1 U4283 ( .A(arr[2099]), .B(n3246), .Y(n7711) );
  OAI21X1 U4284 ( .A(n5509), .B(n3244), .C(n7712), .Y(n10402) );
  NAND2X1 U4285 ( .A(arr[2100]), .B(n3246), .Y(n7712) );
  OAI21X1 U4286 ( .A(n5511), .B(n3245), .C(n7713), .Y(n10403) );
  NAND2X1 U4287 ( .A(arr[2101]), .B(n3246), .Y(n7713) );
  OAI21X1 U4288 ( .A(n5513), .B(n3245), .C(n7714), .Y(n10404) );
  NAND2X1 U4289 ( .A(arr[2102]), .B(n3246), .Y(n7714) );
  OAI21X1 U4290 ( .A(n5515), .B(n3245), .C(n7715), .Y(n10405) );
  NAND2X1 U4291 ( .A(arr[2103]), .B(n3246), .Y(n7715) );
  OAI21X1 U4292 ( .A(n5517), .B(n3244), .C(n7716), .Y(n10406) );
  NAND2X1 U4293 ( .A(arr[2104]), .B(n3247), .Y(n7716) );
  OAI21X1 U4294 ( .A(n5519), .B(n3246), .C(n7717), .Y(n10407) );
  NAND2X1 U4295 ( .A(arr[2105]), .B(n3247), .Y(n7717) );
  OAI21X1 U4296 ( .A(n5521), .B(n3246), .C(n7718), .Y(n10408) );
  NAND2X1 U4297 ( .A(arr[2106]), .B(n3247), .Y(n7718) );
  OAI21X1 U4298 ( .A(n5523), .B(n3245), .C(n7719), .Y(n10409) );
  NAND2X1 U4299 ( .A(arr[2107]), .B(n3247), .Y(n7719) );
  OAI21X1 U4300 ( .A(n5525), .B(n3245), .C(n7720), .Y(n10410) );
  NAND2X1 U4301 ( .A(arr[2108]), .B(n3247), .Y(n7720) );
  OAI21X1 U4302 ( .A(n5527), .B(n3245), .C(n7721), .Y(n10411) );
  NAND2X1 U4303 ( .A(arr[2109]), .B(n3247), .Y(n7721) );
  OAI21X1 U4304 ( .A(n5529), .B(n3245), .C(n7722), .Y(n10412) );
  NAND2X1 U4305 ( .A(arr[2110]), .B(n3247), .Y(n7722) );
  OAI21X1 U4306 ( .A(n5531), .B(n3245), .C(n7723), .Y(n10413) );
  NAND2X1 U4307 ( .A(arr[2111]), .B(n3247), .Y(n7723) );
  OAI21X1 U4308 ( .A(n5533), .B(n3245), .C(n7724), .Y(n10414) );
  NAND2X1 U4309 ( .A(arr[2112]), .B(n3247), .Y(n7724) );
  OAI21X1 U4310 ( .A(n5535), .B(n3245), .C(n7725), .Y(n10415) );
  NAND2X1 U4311 ( .A(arr[2113]), .B(n3247), .Y(n7725) );
  OAI21X1 U4312 ( .A(n5537), .B(n3245), .C(n7726), .Y(n10416) );
  NAND2X1 U4313 ( .A(arr[2114]), .B(n3247), .Y(n7726) );
  OAI21X1 U4314 ( .A(n5539), .B(n3245), .C(n7727), .Y(n10417) );
  NAND2X1 U4315 ( .A(arr[2115]), .B(n3247), .Y(n7727) );
  OAI21X1 U4316 ( .A(n5541), .B(n3245), .C(n7728), .Y(n10418) );
  NAND2X1 U4317 ( .A(arr[2116]), .B(n3247), .Y(n7728) );
  OAI21X1 U4318 ( .A(n5543), .B(n3244), .C(n7729), .Y(n10419) );
  NAND2X1 U4319 ( .A(arr[2117]), .B(n3247), .Y(n7729) );
  OAI21X1 U4320 ( .A(n5545), .B(n3244), .C(n7730), .Y(n10420) );
  NAND2X1 U4321 ( .A(arr[2118]), .B(n3247), .Y(n7730) );
  OAI21X1 U4322 ( .A(n5547), .B(n3244), .C(n7731), .Y(n10421) );
  NAND2X1 U4323 ( .A(arr[2119]), .B(n3247), .Y(n7731) );
  OAI21X1 U4324 ( .A(n5549), .B(n3244), .C(n7732), .Y(n10422) );
  NAND2X1 U4325 ( .A(arr[2120]), .B(n3247), .Y(n7732) );
  OAI21X1 U4326 ( .A(n5551), .B(n3244), .C(n7733), .Y(n10423) );
  NAND2X1 U4327 ( .A(arr[2121]), .B(n3248), .Y(n7733) );
  OAI21X1 U4328 ( .A(n5553), .B(n3244), .C(n7734), .Y(n10424) );
  NAND2X1 U4329 ( .A(arr[2122]), .B(n3248), .Y(n7734) );
  OAI21X1 U4330 ( .A(n5555), .B(n3244), .C(n7735), .Y(n10425) );
  NAND2X1 U4331 ( .A(arr[2123]), .B(n3248), .Y(n7735) );
  OAI21X1 U4332 ( .A(n5557), .B(n3244), .C(n7736), .Y(n10426) );
  NAND2X1 U4333 ( .A(arr[2124]), .B(n3248), .Y(n7736) );
  OAI21X1 U4334 ( .A(n5559), .B(n3243), .C(n7737), .Y(n10427) );
  NAND2X1 U4335 ( .A(arr[2125]), .B(n3248), .Y(n7737) );
  OAI21X1 U4336 ( .A(n5561), .B(n3243), .C(n7738), .Y(n10428) );
  NAND2X1 U4337 ( .A(arr[2126]), .B(n3248), .Y(n7738) );
  OAI21X1 U4338 ( .A(n5563), .B(n3243), .C(n7739), .Y(n10429) );
  NAND2X1 U4339 ( .A(arr[2127]), .B(n3248), .Y(n7739) );
  OAI21X1 U4340 ( .A(n5565), .B(n3243), .C(n7740), .Y(n10430) );
  NAND2X1 U4341 ( .A(arr[2128]), .B(n3248), .Y(n7740) );
  OAI21X1 U4342 ( .A(n5567), .B(n3243), .C(n7741), .Y(n10431) );
  NAND2X1 U4343 ( .A(arr[2129]), .B(n3248), .Y(n7741) );
  OAI21X1 U4344 ( .A(n5569), .B(n3243), .C(n7742), .Y(n10432) );
  NAND2X1 U4345 ( .A(arr[2130]), .B(n3246), .Y(n7742) );
  OAI21X1 U4346 ( .A(n5571), .B(n3243), .C(n7743), .Y(n10433) );
  NAND2X1 U4347 ( .A(arr[2131]), .B(n3246), .Y(n7743) );
  NAND2X1 U4348 ( .A(n7617), .B(n5703), .Y(n7702) );
  NOR2X1 U4350 ( .A(wr_ptr[2]), .B(wr_ptr[3]), .Y(n5705) );
  OAI21X1 U4351 ( .A(n5491), .B(n3237), .C(n7746), .Y(n10434) );
  NAND2X1 U4352 ( .A(arr[2132]), .B(n3240), .Y(n7746) );
  OAI21X1 U4353 ( .A(n5493), .B(n3237), .C(n7747), .Y(n10435) );
  NAND2X1 U4354 ( .A(arr[2133]), .B(n3240), .Y(n7747) );
  OAI21X1 U4355 ( .A(n5495), .B(n3237), .C(n7748), .Y(n10436) );
  NAND2X1 U4356 ( .A(arr[2134]), .B(n3240), .Y(n7748) );
  OAI21X1 U4357 ( .A(n5497), .B(n3237), .C(n7749), .Y(n10437) );
  NAND2X1 U4358 ( .A(arr[2135]), .B(n3240), .Y(n7749) );
  OAI21X1 U4359 ( .A(n5499), .B(n3237), .C(n7750), .Y(n10438) );
  NAND2X1 U4360 ( .A(arr[2136]), .B(n3240), .Y(n7750) );
  OAI21X1 U4361 ( .A(n5501), .B(n3238), .C(n7751), .Y(n10439) );
  NAND2X1 U4362 ( .A(arr[2137]), .B(n3240), .Y(n7751) );
  OAI21X1 U4363 ( .A(n5503), .B(n3238), .C(n7752), .Y(n10440) );
  NAND2X1 U4364 ( .A(arr[2138]), .B(n3240), .Y(n7752) );
  OAI21X1 U4365 ( .A(n5505), .B(n3238), .C(n7753), .Y(n10441) );
  NAND2X1 U4366 ( .A(arr[2139]), .B(n3240), .Y(n7753) );
  OAI21X1 U4367 ( .A(n5507), .B(n3237), .C(n7754), .Y(n10442) );
  NAND2X1 U4368 ( .A(arr[2140]), .B(n3240), .Y(n7754) );
  OAI21X1 U4369 ( .A(n5509), .B(n3238), .C(n7755), .Y(n10443) );
  NAND2X1 U4370 ( .A(arr[2141]), .B(n3240), .Y(n7755) );
  OAI21X1 U4371 ( .A(n5511), .B(n3239), .C(n7756), .Y(n10444) );
  NAND2X1 U4372 ( .A(arr[2142]), .B(n3240), .Y(n7756) );
  OAI21X1 U4373 ( .A(n5513), .B(n3239), .C(n7757), .Y(n10445) );
  NAND2X1 U4374 ( .A(arr[2143]), .B(n3240), .Y(n7757) );
  OAI21X1 U4375 ( .A(n5515), .B(n3239), .C(n7758), .Y(n10446) );
  NAND2X1 U4376 ( .A(arr[2144]), .B(n3240), .Y(n7758) );
  OAI21X1 U4377 ( .A(n5517), .B(n3238), .C(n7759), .Y(n10447) );
  NAND2X1 U4378 ( .A(arr[2145]), .B(n3241), .Y(n7759) );
  OAI21X1 U4379 ( .A(n5519), .B(n3240), .C(n7760), .Y(n10448) );
  NAND2X1 U4380 ( .A(arr[2146]), .B(n3241), .Y(n7760) );
  OAI21X1 U4381 ( .A(n5521), .B(n3240), .C(n7761), .Y(n10449) );
  NAND2X1 U4382 ( .A(arr[2147]), .B(n3241), .Y(n7761) );
  OAI21X1 U4383 ( .A(n5523), .B(n3239), .C(n7762), .Y(n10450) );
  NAND2X1 U4384 ( .A(arr[2148]), .B(n3241), .Y(n7762) );
  OAI21X1 U4385 ( .A(n5525), .B(n3239), .C(n7763), .Y(n10451) );
  NAND2X1 U4386 ( .A(arr[2149]), .B(n3241), .Y(n7763) );
  OAI21X1 U4387 ( .A(n5527), .B(n3239), .C(n7764), .Y(n10452) );
  NAND2X1 U4388 ( .A(arr[2150]), .B(n3241), .Y(n7764) );
  OAI21X1 U4389 ( .A(n5529), .B(n3239), .C(n7765), .Y(n10453) );
  NAND2X1 U4390 ( .A(arr[2151]), .B(n3241), .Y(n7765) );
  OAI21X1 U4391 ( .A(n5531), .B(n3239), .C(n7766), .Y(n10454) );
  NAND2X1 U4392 ( .A(arr[2152]), .B(n3241), .Y(n7766) );
  OAI21X1 U4393 ( .A(n5533), .B(n3239), .C(n7767), .Y(n10455) );
  NAND2X1 U4394 ( .A(arr[2153]), .B(n3241), .Y(n7767) );
  OAI21X1 U4395 ( .A(n5535), .B(n3239), .C(n7768), .Y(n10456) );
  NAND2X1 U4396 ( .A(arr[2154]), .B(n3241), .Y(n7768) );
  OAI21X1 U4397 ( .A(n5537), .B(n3239), .C(n7769), .Y(n10457) );
  NAND2X1 U4398 ( .A(arr[2155]), .B(n3241), .Y(n7769) );
  OAI21X1 U4399 ( .A(n5539), .B(n3239), .C(n7770), .Y(n10458) );
  NAND2X1 U4400 ( .A(arr[2156]), .B(n3241), .Y(n7770) );
  OAI21X1 U4401 ( .A(n5541), .B(n3239), .C(n7771), .Y(n10459) );
  NAND2X1 U4402 ( .A(arr[2157]), .B(n3241), .Y(n7771) );
  OAI21X1 U4403 ( .A(n5543), .B(n3238), .C(n7772), .Y(n10460) );
  NAND2X1 U4404 ( .A(arr[2158]), .B(n3241), .Y(n7772) );
  OAI21X1 U4405 ( .A(n5545), .B(n3238), .C(n7773), .Y(n10461) );
  NAND2X1 U4406 ( .A(arr[2159]), .B(n3241), .Y(n7773) );
  OAI21X1 U4407 ( .A(n5547), .B(n3238), .C(n7774), .Y(n10462) );
  NAND2X1 U4408 ( .A(arr[2160]), .B(n3241), .Y(n7774) );
  OAI21X1 U4409 ( .A(n5549), .B(n3238), .C(n7775), .Y(n10463) );
  NAND2X1 U4410 ( .A(arr[2161]), .B(n3241), .Y(n7775) );
  OAI21X1 U4411 ( .A(n5551), .B(n3238), .C(n7776), .Y(n10464) );
  NAND2X1 U4412 ( .A(arr[2162]), .B(n3242), .Y(n7776) );
  OAI21X1 U4413 ( .A(n5553), .B(n3238), .C(n7777), .Y(n10465) );
  NAND2X1 U4414 ( .A(arr[2163]), .B(n3242), .Y(n7777) );
  OAI21X1 U4415 ( .A(n5555), .B(n3238), .C(n7778), .Y(n10466) );
  NAND2X1 U4416 ( .A(arr[2164]), .B(n3242), .Y(n7778) );
  OAI21X1 U4417 ( .A(n5557), .B(n3238), .C(n7779), .Y(n10467) );
  NAND2X1 U4418 ( .A(arr[2165]), .B(n3242), .Y(n7779) );
  OAI21X1 U4419 ( .A(n5559), .B(n3237), .C(n7780), .Y(n10468) );
  NAND2X1 U4420 ( .A(arr[2166]), .B(n3242), .Y(n7780) );
  OAI21X1 U4421 ( .A(n5561), .B(n3237), .C(n7781), .Y(n10469) );
  NAND2X1 U4422 ( .A(arr[2167]), .B(n3242), .Y(n7781) );
  OAI21X1 U4423 ( .A(n5563), .B(n3237), .C(n7782), .Y(n10470) );
  NAND2X1 U4424 ( .A(arr[2168]), .B(n3242), .Y(n7782) );
  OAI21X1 U4425 ( .A(n5565), .B(n3237), .C(n7783), .Y(n10471) );
  NAND2X1 U4426 ( .A(arr[2169]), .B(n3242), .Y(n7783) );
  OAI21X1 U4427 ( .A(n5567), .B(n3237), .C(n7784), .Y(n10472) );
  NAND2X1 U4428 ( .A(arr[2170]), .B(n3242), .Y(n7784) );
  OAI21X1 U4429 ( .A(n5569), .B(n3237), .C(n7785), .Y(n10473) );
  NAND2X1 U4430 ( .A(arr[2171]), .B(n3240), .Y(n7785) );
  OAI21X1 U4431 ( .A(n5571), .B(n3237), .C(n7786), .Y(n10474) );
  NAND2X1 U4432 ( .A(arr[2172]), .B(n3240), .Y(n7786) );
  NAND2X1 U4433 ( .A(n7787), .B(n5573), .Y(n7745) );
  OAI21X1 U4434 ( .A(n5491), .B(n3231), .C(n7789), .Y(n10475) );
  NAND2X1 U4435 ( .A(arr[2173]), .B(n3234), .Y(n7789) );
  OAI21X1 U4436 ( .A(n5493), .B(n3231), .C(n7790), .Y(n10476) );
  NAND2X1 U4437 ( .A(arr[2174]), .B(n3234), .Y(n7790) );
  OAI21X1 U4438 ( .A(n5495), .B(n3231), .C(n7791), .Y(n10477) );
  NAND2X1 U4439 ( .A(arr[2175]), .B(n3234), .Y(n7791) );
  OAI21X1 U4440 ( .A(n5497), .B(n3231), .C(n7792), .Y(n10478) );
  NAND2X1 U4441 ( .A(arr[2176]), .B(n3234), .Y(n7792) );
  OAI21X1 U4442 ( .A(n5499), .B(n3231), .C(n7793), .Y(n10479) );
  NAND2X1 U4443 ( .A(arr[2177]), .B(n3234), .Y(n7793) );
  OAI21X1 U4444 ( .A(n5501), .B(n3232), .C(n7794), .Y(n10480) );
  NAND2X1 U4445 ( .A(arr[2178]), .B(n3234), .Y(n7794) );
  OAI21X1 U4446 ( .A(n5503), .B(n3232), .C(n7795), .Y(n10481) );
  NAND2X1 U4447 ( .A(arr[2179]), .B(n3234), .Y(n7795) );
  OAI21X1 U4448 ( .A(n5505), .B(n3232), .C(n7796), .Y(n10482) );
  NAND2X1 U4449 ( .A(arr[2180]), .B(n3234), .Y(n7796) );
  OAI21X1 U4450 ( .A(n5507), .B(n3231), .C(n7797), .Y(n10483) );
  NAND2X1 U4451 ( .A(arr[2181]), .B(n3234), .Y(n7797) );
  OAI21X1 U4452 ( .A(n5509), .B(n3232), .C(n7798), .Y(n10484) );
  NAND2X1 U4453 ( .A(arr[2182]), .B(n3234), .Y(n7798) );
  OAI21X1 U4454 ( .A(n5511), .B(n3233), .C(n7799), .Y(n10485) );
  NAND2X1 U4455 ( .A(arr[2183]), .B(n3234), .Y(n7799) );
  OAI21X1 U4456 ( .A(n5513), .B(n3233), .C(n7800), .Y(n10486) );
  NAND2X1 U4457 ( .A(arr[2184]), .B(n3234), .Y(n7800) );
  OAI21X1 U4458 ( .A(n5515), .B(n3233), .C(n7801), .Y(n10487) );
  NAND2X1 U4459 ( .A(arr[2185]), .B(n3234), .Y(n7801) );
  OAI21X1 U4460 ( .A(n5517), .B(n3232), .C(n7802), .Y(n10488) );
  NAND2X1 U4461 ( .A(arr[2186]), .B(n3235), .Y(n7802) );
  OAI21X1 U4462 ( .A(n5519), .B(n3234), .C(n7803), .Y(n10489) );
  NAND2X1 U4463 ( .A(arr[2187]), .B(n3235), .Y(n7803) );
  OAI21X1 U4464 ( .A(n5521), .B(n3234), .C(n7804), .Y(n10490) );
  NAND2X1 U4465 ( .A(arr[2188]), .B(n3235), .Y(n7804) );
  OAI21X1 U4466 ( .A(n5523), .B(n3233), .C(n7805), .Y(n10491) );
  NAND2X1 U4467 ( .A(arr[2189]), .B(n3235), .Y(n7805) );
  OAI21X1 U4468 ( .A(n5525), .B(n3233), .C(n7806), .Y(n10492) );
  NAND2X1 U4469 ( .A(arr[2190]), .B(n3235), .Y(n7806) );
  OAI21X1 U4470 ( .A(n5527), .B(n3233), .C(n7807), .Y(n10493) );
  NAND2X1 U4471 ( .A(arr[2191]), .B(n3235), .Y(n7807) );
  OAI21X1 U4472 ( .A(n5529), .B(n3233), .C(n7808), .Y(n10494) );
  NAND2X1 U4473 ( .A(arr[2192]), .B(n3235), .Y(n7808) );
  OAI21X1 U4474 ( .A(n5531), .B(n3233), .C(n7809), .Y(n10495) );
  NAND2X1 U4475 ( .A(arr[2193]), .B(n3235), .Y(n7809) );
  OAI21X1 U4476 ( .A(n5533), .B(n3233), .C(n7810), .Y(n10496) );
  NAND2X1 U4477 ( .A(arr[2194]), .B(n3235), .Y(n7810) );
  OAI21X1 U4478 ( .A(n5535), .B(n3233), .C(n7811), .Y(n10497) );
  NAND2X1 U4479 ( .A(arr[2195]), .B(n3235), .Y(n7811) );
  OAI21X1 U4480 ( .A(n5537), .B(n3233), .C(n7812), .Y(n10498) );
  NAND2X1 U4481 ( .A(arr[2196]), .B(n3235), .Y(n7812) );
  OAI21X1 U4482 ( .A(n5539), .B(n3233), .C(n7813), .Y(n10499) );
  NAND2X1 U4483 ( .A(arr[2197]), .B(n3235), .Y(n7813) );
  OAI21X1 U4484 ( .A(n5541), .B(n3233), .C(n7814), .Y(n10500) );
  NAND2X1 U4485 ( .A(arr[2198]), .B(n3235), .Y(n7814) );
  OAI21X1 U4486 ( .A(n5543), .B(n3232), .C(n7815), .Y(n10501) );
  NAND2X1 U4487 ( .A(arr[2199]), .B(n3235), .Y(n7815) );
  OAI21X1 U4488 ( .A(n5545), .B(n3232), .C(n7816), .Y(n10502) );
  NAND2X1 U4489 ( .A(arr[2200]), .B(n3235), .Y(n7816) );
  OAI21X1 U4490 ( .A(n5547), .B(n3232), .C(n7817), .Y(n10503) );
  NAND2X1 U4491 ( .A(arr[2201]), .B(n3235), .Y(n7817) );
  OAI21X1 U4492 ( .A(n5549), .B(n3232), .C(n7818), .Y(n10504) );
  NAND2X1 U4493 ( .A(arr[2202]), .B(n3235), .Y(n7818) );
  OAI21X1 U4494 ( .A(n5551), .B(n3232), .C(n7819), .Y(n10505) );
  NAND2X1 U4495 ( .A(arr[2203]), .B(n3236), .Y(n7819) );
  OAI21X1 U4496 ( .A(n5553), .B(n3232), .C(n7820), .Y(n10506) );
  NAND2X1 U4497 ( .A(arr[2204]), .B(n3236), .Y(n7820) );
  OAI21X1 U4498 ( .A(n5555), .B(n3232), .C(n7821), .Y(n10507) );
  NAND2X1 U4499 ( .A(arr[2205]), .B(n3236), .Y(n7821) );
  OAI21X1 U4500 ( .A(n5557), .B(n3232), .C(n7822), .Y(n10508) );
  NAND2X1 U4501 ( .A(arr[2206]), .B(n3236), .Y(n7822) );
  OAI21X1 U4502 ( .A(n5559), .B(n3231), .C(n7823), .Y(n10509) );
  NAND2X1 U4503 ( .A(arr[2207]), .B(n3236), .Y(n7823) );
  OAI21X1 U4504 ( .A(n5561), .B(n3231), .C(n7824), .Y(n10510) );
  NAND2X1 U4505 ( .A(arr[2208]), .B(n3236), .Y(n7824) );
  OAI21X1 U4506 ( .A(n5563), .B(n3231), .C(n7825), .Y(n10511) );
  NAND2X1 U4507 ( .A(arr[2209]), .B(n3236), .Y(n7825) );
  OAI21X1 U4508 ( .A(n5565), .B(n3231), .C(n7826), .Y(n10512) );
  NAND2X1 U4509 ( .A(arr[2210]), .B(n3236), .Y(n7826) );
  OAI21X1 U4510 ( .A(n5567), .B(n3231), .C(n7827), .Y(n10513) );
  NAND2X1 U4511 ( .A(arr[2211]), .B(n3236), .Y(n7827) );
  OAI21X1 U4512 ( .A(n5569), .B(n3231), .C(n7828), .Y(n10514) );
  NAND2X1 U4513 ( .A(arr[2212]), .B(n3234), .Y(n7828) );
  OAI21X1 U4514 ( .A(n5571), .B(n3231), .C(n7829), .Y(n10515) );
  NAND2X1 U4515 ( .A(arr[2213]), .B(n3234), .Y(n7829) );
  NAND2X1 U4516 ( .A(n7787), .B(n5617), .Y(n7788) );
  OAI21X1 U4517 ( .A(n5491), .B(n3225), .C(n7831), .Y(n10516) );
  NAND2X1 U4518 ( .A(arr[2214]), .B(n3228), .Y(n7831) );
  OAI21X1 U4519 ( .A(n5493), .B(n3225), .C(n7832), .Y(n10517) );
  NAND2X1 U4520 ( .A(arr[2215]), .B(n3228), .Y(n7832) );
  OAI21X1 U4521 ( .A(n5495), .B(n3225), .C(n7833), .Y(n10518) );
  NAND2X1 U4522 ( .A(arr[2216]), .B(n3228), .Y(n7833) );
  OAI21X1 U4523 ( .A(n5497), .B(n3225), .C(n7834), .Y(n10519) );
  NAND2X1 U4524 ( .A(arr[2217]), .B(n3228), .Y(n7834) );
  OAI21X1 U4525 ( .A(n5499), .B(n3225), .C(n7835), .Y(n10520) );
  NAND2X1 U4526 ( .A(arr[2218]), .B(n3228), .Y(n7835) );
  OAI21X1 U4527 ( .A(n5501), .B(n3226), .C(n7836), .Y(n10521) );
  NAND2X1 U4528 ( .A(arr[2219]), .B(n3228), .Y(n7836) );
  OAI21X1 U4529 ( .A(n5503), .B(n3226), .C(n7837), .Y(n10522) );
  NAND2X1 U4530 ( .A(arr[2220]), .B(n3228), .Y(n7837) );
  OAI21X1 U4531 ( .A(n5505), .B(n3226), .C(n7838), .Y(n10523) );
  NAND2X1 U4532 ( .A(arr[2221]), .B(n3228), .Y(n7838) );
  OAI21X1 U4533 ( .A(n5507), .B(n3225), .C(n7839), .Y(n10524) );
  NAND2X1 U4534 ( .A(arr[2222]), .B(n3228), .Y(n7839) );
  OAI21X1 U4535 ( .A(n5509), .B(n3226), .C(n7840), .Y(n10525) );
  NAND2X1 U4536 ( .A(arr[2223]), .B(n3228), .Y(n7840) );
  OAI21X1 U4537 ( .A(n5511), .B(n3227), .C(n7841), .Y(n10526) );
  NAND2X1 U4538 ( .A(arr[2224]), .B(n3228), .Y(n7841) );
  OAI21X1 U4539 ( .A(n5513), .B(n3227), .C(n7842), .Y(n10527) );
  NAND2X1 U4540 ( .A(arr[2225]), .B(n3228), .Y(n7842) );
  OAI21X1 U4541 ( .A(n5515), .B(n3227), .C(n7843), .Y(n10528) );
  NAND2X1 U4542 ( .A(arr[2226]), .B(n3228), .Y(n7843) );
  OAI21X1 U4543 ( .A(n5517), .B(n3226), .C(n7844), .Y(n10529) );
  NAND2X1 U4544 ( .A(arr[2227]), .B(n3229), .Y(n7844) );
  OAI21X1 U4545 ( .A(n5519), .B(n3228), .C(n7845), .Y(n10530) );
  NAND2X1 U4546 ( .A(arr[2228]), .B(n3229), .Y(n7845) );
  OAI21X1 U4547 ( .A(n5521), .B(n3228), .C(n7846), .Y(n10531) );
  NAND2X1 U4548 ( .A(arr[2229]), .B(n3229), .Y(n7846) );
  OAI21X1 U4549 ( .A(n5523), .B(n3227), .C(n7847), .Y(n10532) );
  NAND2X1 U4550 ( .A(arr[2230]), .B(n3229), .Y(n7847) );
  OAI21X1 U4551 ( .A(n5525), .B(n3227), .C(n7848), .Y(n10533) );
  NAND2X1 U4552 ( .A(arr[2231]), .B(n3229), .Y(n7848) );
  OAI21X1 U4553 ( .A(n5527), .B(n3227), .C(n7849), .Y(n10534) );
  NAND2X1 U4554 ( .A(arr[2232]), .B(n3229), .Y(n7849) );
  OAI21X1 U4555 ( .A(n5529), .B(n3227), .C(n7850), .Y(n10535) );
  NAND2X1 U4556 ( .A(arr[2233]), .B(n3229), .Y(n7850) );
  OAI21X1 U4557 ( .A(n5531), .B(n3227), .C(n7851), .Y(n10536) );
  NAND2X1 U4558 ( .A(arr[2234]), .B(n3229), .Y(n7851) );
  OAI21X1 U4559 ( .A(n5533), .B(n3227), .C(n7852), .Y(n10537) );
  NAND2X1 U4560 ( .A(arr[2235]), .B(n3229), .Y(n7852) );
  OAI21X1 U4561 ( .A(n5535), .B(n3227), .C(n7853), .Y(n10538) );
  NAND2X1 U4562 ( .A(arr[2236]), .B(n3229), .Y(n7853) );
  OAI21X1 U4563 ( .A(n5537), .B(n3227), .C(n7854), .Y(n10539) );
  NAND2X1 U4564 ( .A(arr[2237]), .B(n3229), .Y(n7854) );
  OAI21X1 U4565 ( .A(n5539), .B(n3227), .C(n7855), .Y(n10540) );
  NAND2X1 U4566 ( .A(arr[2238]), .B(n3229), .Y(n7855) );
  OAI21X1 U4567 ( .A(n5541), .B(n3227), .C(n7856), .Y(n10541) );
  NAND2X1 U4568 ( .A(arr[2239]), .B(n3229), .Y(n7856) );
  OAI21X1 U4569 ( .A(n5543), .B(n3226), .C(n7857), .Y(n10542) );
  NAND2X1 U4570 ( .A(arr[2240]), .B(n3229), .Y(n7857) );
  OAI21X1 U4571 ( .A(n5545), .B(n3226), .C(n7858), .Y(n10543) );
  NAND2X1 U4572 ( .A(arr[2241]), .B(n3229), .Y(n7858) );
  OAI21X1 U4573 ( .A(n5547), .B(n3226), .C(n7859), .Y(n10544) );
  NAND2X1 U4574 ( .A(arr[2242]), .B(n3229), .Y(n7859) );
  OAI21X1 U4575 ( .A(n5549), .B(n3226), .C(n7860), .Y(n10545) );
  NAND2X1 U4576 ( .A(arr[2243]), .B(n3229), .Y(n7860) );
  OAI21X1 U4577 ( .A(n5551), .B(n3226), .C(n7861), .Y(n10546) );
  NAND2X1 U4578 ( .A(arr[2244]), .B(n3230), .Y(n7861) );
  OAI21X1 U4579 ( .A(n5553), .B(n3226), .C(n7862), .Y(n10547) );
  NAND2X1 U4580 ( .A(arr[2245]), .B(n3230), .Y(n7862) );
  OAI21X1 U4581 ( .A(n5555), .B(n3226), .C(n7863), .Y(n10548) );
  NAND2X1 U4582 ( .A(arr[2246]), .B(n3230), .Y(n7863) );
  OAI21X1 U4583 ( .A(n5557), .B(n3226), .C(n7864), .Y(n10549) );
  NAND2X1 U4584 ( .A(arr[2247]), .B(n3230), .Y(n7864) );
  OAI21X1 U4585 ( .A(n5559), .B(n3225), .C(n7865), .Y(n10550) );
  NAND2X1 U4586 ( .A(arr[2248]), .B(n3230), .Y(n7865) );
  OAI21X1 U4587 ( .A(n5561), .B(n3225), .C(n7866), .Y(n10551) );
  NAND2X1 U4588 ( .A(arr[2249]), .B(n3230), .Y(n7866) );
  OAI21X1 U4589 ( .A(n5563), .B(n3225), .C(n7867), .Y(n10552) );
  NAND2X1 U4590 ( .A(arr[2250]), .B(n3230), .Y(n7867) );
  OAI21X1 U4591 ( .A(n5565), .B(n3225), .C(n7868), .Y(n10553) );
  NAND2X1 U4592 ( .A(arr[2251]), .B(n3230), .Y(n7868) );
  OAI21X1 U4593 ( .A(n5567), .B(n3225), .C(n7869), .Y(n10554) );
  NAND2X1 U4594 ( .A(arr[2252]), .B(n3230), .Y(n7869) );
  OAI21X1 U4595 ( .A(n5569), .B(n3225), .C(n7870), .Y(n10555) );
  NAND2X1 U4596 ( .A(arr[2253]), .B(n3228), .Y(n7870) );
  OAI21X1 U4597 ( .A(n5571), .B(n3225), .C(n7871), .Y(n10556) );
  NAND2X1 U4598 ( .A(arr[2254]), .B(n3228), .Y(n7871) );
  NAND2X1 U4599 ( .A(n7787), .B(n5660), .Y(n7830) );
  OAI21X1 U4600 ( .A(n5491), .B(n3219), .C(n7873), .Y(n10557) );
  NAND2X1 U4601 ( .A(arr[2255]), .B(n3222), .Y(n7873) );
  OAI21X1 U4602 ( .A(n5493), .B(n3219), .C(n7874), .Y(n10558) );
  NAND2X1 U4603 ( .A(arr[2256]), .B(n3222), .Y(n7874) );
  OAI21X1 U4604 ( .A(n5495), .B(n3219), .C(n7875), .Y(n10559) );
  NAND2X1 U4605 ( .A(arr[2257]), .B(n3222), .Y(n7875) );
  OAI21X1 U4606 ( .A(n5497), .B(n3219), .C(n7876), .Y(n10560) );
  NAND2X1 U4607 ( .A(arr[2258]), .B(n3222), .Y(n7876) );
  OAI21X1 U4608 ( .A(n5499), .B(n3219), .C(n7877), .Y(n10561) );
  NAND2X1 U4609 ( .A(arr[2259]), .B(n3222), .Y(n7877) );
  OAI21X1 U4610 ( .A(n5501), .B(n3220), .C(n7878), .Y(n10562) );
  NAND2X1 U4611 ( .A(arr[2260]), .B(n3222), .Y(n7878) );
  OAI21X1 U4612 ( .A(n5503), .B(n3220), .C(n7879), .Y(n10563) );
  NAND2X1 U4613 ( .A(arr[2261]), .B(n3222), .Y(n7879) );
  OAI21X1 U4614 ( .A(n5505), .B(n3220), .C(n7880), .Y(n10564) );
  NAND2X1 U4615 ( .A(arr[2262]), .B(n3222), .Y(n7880) );
  OAI21X1 U4616 ( .A(n5507), .B(n3219), .C(n7881), .Y(n10565) );
  NAND2X1 U4617 ( .A(arr[2263]), .B(n3222), .Y(n7881) );
  OAI21X1 U4618 ( .A(n5509), .B(n3220), .C(n7882), .Y(n10566) );
  NAND2X1 U4619 ( .A(arr[2264]), .B(n3222), .Y(n7882) );
  OAI21X1 U4620 ( .A(n5511), .B(n3221), .C(n7883), .Y(n10567) );
  NAND2X1 U4621 ( .A(arr[2265]), .B(n3222), .Y(n7883) );
  OAI21X1 U4622 ( .A(n5513), .B(n3221), .C(n7884), .Y(n10568) );
  NAND2X1 U4623 ( .A(arr[2266]), .B(n3222), .Y(n7884) );
  OAI21X1 U4624 ( .A(n5515), .B(n3221), .C(n7885), .Y(n10569) );
  NAND2X1 U4625 ( .A(arr[2267]), .B(n3222), .Y(n7885) );
  OAI21X1 U4626 ( .A(n5517), .B(n3220), .C(n7886), .Y(n10570) );
  NAND2X1 U4627 ( .A(arr[2268]), .B(n3223), .Y(n7886) );
  OAI21X1 U4628 ( .A(n5519), .B(n3222), .C(n7887), .Y(n10571) );
  NAND2X1 U4629 ( .A(arr[2269]), .B(n3223), .Y(n7887) );
  OAI21X1 U4630 ( .A(n5521), .B(n3222), .C(n7888), .Y(n10572) );
  NAND2X1 U4631 ( .A(arr[2270]), .B(n3223), .Y(n7888) );
  OAI21X1 U4632 ( .A(n5523), .B(n3221), .C(n7889), .Y(n10573) );
  NAND2X1 U4633 ( .A(arr[2271]), .B(n3223), .Y(n7889) );
  OAI21X1 U4634 ( .A(n5525), .B(n3221), .C(n7890), .Y(n10574) );
  NAND2X1 U4635 ( .A(arr[2272]), .B(n3223), .Y(n7890) );
  OAI21X1 U4636 ( .A(n5527), .B(n3221), .C(n7891), .Y(n10575) );
  NAND2X1 U4637 ( .A(arr[2273]), .B(n3223), .Y(n7891) );
  OAI21X1 U4638 ( .A(n5529), .B(n3221), .C(n7892), .Y(n10576) );
  NAND2X1 U4639 ( .A(arr[2274]), .B(n3223), .Y(n7892) );
  OAI21X1 U4640 ( .A(n5531), .B(n3221), .C(n7893), .Y(n10577) );
  NAND2X1 U4641 ( .A(arr[2275]), .B(n3223), .Y(n7893) );
  OAI21X1 U4642 ( .A(n5533), .B(n3221), .C(n7894), .Y(n10578) );
  NAND2X1 U4643 ( .A(arr[2276]), .B(n3223), .Y(n7894) );
  OAI21X1 U4644 ( .A(n5535), .B(n3221), .C(n7895), .Y(n10579) );
  NAND2X1 U4645 ( .A(arr[2277]), .B(n3223), .Y(n7895) );
  OAI21X1 U4646 ( .A(n5537), .B(n3221), .C(n7896), .Y(n10580) );
  NAND2X1 U4647 ( .A(arr[2278]), .B(n3223), .Y(n7896) );
  OAI21X1 U4648 ( .A(n5539), .B(n3221), .C(n7897), .Y(n10581) );
  NAND2X1 U4649 ( .A(arr[2279]), .B(n3223), .Y(n7897) );
  OAI21X1 U4650 ( .A(n5541), .B(n3221), .C(n7898), .Y(n10582) );
  NAND2X1 U4651 ( .A(arr[2280]), .B(n3223), .Y(n7898) );
  OAI21X1 U4652 ( .A(n5543), .B(n3220), .C(n7899), .Y(n10583) );
  NAND2X1 U4653 ( .A(arr[2281]), .B(n3223), .Y(n7899) );
  OAI21X1 U4654 ( .A(n5545), .B(n3220), .C(n7900), .Y(n10584) );
  NAND2X1 U4655 ( .A(arr[2282]), .B(n3223), .Y(n7900) );
  OAI21X1 U4656 ( .A(n5547), .B(n3220), .C(n7901), .Y(n10585) );
  NAND2X1 U4657 ( .A(arr[2283]), .B(n3223), .Y(n7901) );
  OAI21X1 U4658 ( .A(n5549), .B(n3220), .C(n7902), .Y(n10586) );
  NAND2X1 U4659 ( .A(arr[2284]), .B(n3223), .Y(n7902) );
  OAI21X1 U4660 ( .A(n5551), .B(n3220), .C(n7903), .Y(n10587) );
  NAND2X1 U4661 ( .A(arr[2285]), .B(n3224), .Y(n7903) );
  OAI21X1 U4662 ( .A(n5553), .B(n3220), .C(n7904), .Y(n10588) );
  NAND2X1 U4663 ( .A(arr[2286]), .B(n3224), .Y(n7904) );
  OAI21X1 U4664 ( .A(n5555), .B(n3220), .C(n7905), .Y(n10589) );
  NAND2X1 U4665 ( .A(arr[2287]), .B(n3224), .Y(n7905) );
  OAI21X1 U4666 ( .A(n5557), .B(n3220), .C(n7906), .Y(n10590) );
  NAND2X1 U4667 ( .A(arr[2288]), .B(n3224), .Y(n7906) );
  OAI21X1 U4668 ( .A(n5559), .B(n3219), .C(n7907), .Y(n10591) );
  NAND2X1 U4669 ( .A(arr[2289]), .B(n3224), .Y(n7907) );
  OAI21X1 U4670 ( .A(n5561), .B(n3219), .C(n7908), .Y(n10592) );
  NAND2X1 U4671 ( .A(arr[2290]), .B(n3224), .Y(n7908) );
  OAI21X1 U4672 ( .A(n5563), .B(n3219), .C(n7909), .Y(n10593) );
  NAND2X1 U4673 ( .A(arr[2291]), .B(n3224), .Y(n7909) );
  OAI21X1 U4674 ( .A(n5565), .B(n3219), .C(n7910), .Y(n10594) );
  NAND2X1 U4675 ( .A(arr[2292]), .B(n3224), .Y(n7910) );
  OAI21X1 U4676 ( .A(n5567), .B(n3219), .C(n7911), .Y(n10595) );
  NAND2X1 U4677 ( .A(arr[2293]), .B(n3224), .Y(n7911) );
  OAI21X1 U4678 ( .A(n5569), .B(n3219), .C(n7912), .Y(n10596) );
  NAND2X1 U4679 ( .A(arr[2294]), .B(n3222), .Y(n7912) );
  OAI21X1 U4680 ( .A(n5571), .B(n3219), .C(n7913), .Y(n10597) );
  NAND2X1 U4681 ( .A(arr[2295]), .B(n3222), .Y(n7913) );
  NAND2X1 U4682 ( .A(n7787), .B(n5703), .Y(n7872) );
  NOR2X1 U4684 ( .A(n7914), .B(wr_ptr[3]), .Y(n5875) );
  OAI21X1 U4763 ( .A(n5569), .B(n3215), .C(n7955), .Y(n10637) );
  NAND2X1 U4764 ( .A(arr[2335]), .B(n3216), .Y(n7955) );
  OAI21X1 U4765 ( .A(n5571), .B(n3215), .C(n7956), .Y(n10638) );
  NAND2X1 U4766 ( .A(arr[2336]), .B(n3216), .Y(n7956) );
  NAND2X1 U4767 ( .A(n7957), .B(n5573), .Y(n7915) );
  OAI21X1 U4846 ( .A(n5569), .B(n3211), .C(n7998), .Y(n10678) );
  NAND2X1 U4847 ( .A(arr[2376]), .B(n3212), .Y(n7998) );
  OAI21X1 U4848 ( .A(n5571), .B(n3211), .C(n7999), .Y(n10679) );
  NAND2X1 U4849 ( .A(arr[2377]), .B(n3212), .Y(n7999) );
  NAND2X1 U4850 ( .A(n7957), .B(n5617), .Y(n7958) );
  OAI21X1 U4929 ( .A(n5569), .B(n3207), .C(n8040), .Y(n10719) );
  NAND2X1 U4930 ( .A(arr[2417]), .B(n3208), .Y(n8040) );
  OAI21X1 U4931 ( .A(n5571), .B(n3207), .C(n8041), .Y(n10720) );
  NAND2X1 U4932 ( .A(arr[2418]), .B(n3208), .Y(n8041) );
  NAND2X1 U4933 ( .A(n7957), .B(n5660), .Y(n8000) );
  OAI21X1 U5012 ( .A(n5569), .B(n3203), .C(n8082), .Y(n10760) );
  NAND2X1 U5013 ( .A(arr[2458]), .B(n3204), .Y(n8082) );
  OAI21X1 U5014 ( .A(n5571), .B(n3203), .C(n8083), .Y(n10761) );
  NAND2X1 U5015 ( .A(arr[2459]), .B(n3204), .Y(n8083) );
  NAND2X1 U5016 ( .A(n7957), .B(n5703), .Y(n8042) );
  NOR2X1 U5018 ( .A(n8084), .B(wr_ptr[2]), .Y(n6045) );
  OAI21X1 U5097 ( .A(n5569), .B(n3199), .C(n8125), .Y(n10801) );
  NAND2X1 U5098 ( .A(arr[2499]), .B(n3200), .Y(n8125) );
  OAI21X1 U5099 ( .A(n5571), .B(n3199), .C(n8126), .Y(n10802) );
  NAND2X1 U5100 ( .A(arr[2500]), .B(n3200), .Y(n8126) );
  NAND2X1 U5101 ( .A(n8127), .B(n5573), .Y(n8085) );
  NOR2X1 U5102 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .Y(n5573) );
  OAI21X1 U5181 ( .A(n5569), .B(n3195), .C(n8168), .Y(n10842) );
  NAND2X1 U5182 ( .A(arr[2540]), .B(n3196), .Y(n8168) );
  OAI21X1 U5183 ( .A(n5571), .B(n3195), .C(n8169), .Y(n10843) );
  NAND2X1 U5184 ( .A(arr[2541]), .B(n3196), .Y(n8169) );
  NAND2X1 U5185 ( .A(n8127), .B(n5617), .Y(n8128) );
  NOR2X1 U5186 ( .A(n8170), .B(wr_ptr[1]), .Y(n5617) );
  OAI21X1 U5265 ( .A(n5569), .B(n3191), .C(n8211), .Y(n10883) );
  NAND2X1 U5266 ( .A(arr[2581]), .B(n3192), .Y(n8211) );
  OAI21X1 U5267 ( .A(n5571), .B(n3191), .C(n8212), .Y(n10884) );
  NAND2X1 U5268 ( .A(arr[2582]), .B(n3192), .Y(n8212) );
  NAND2X1 U5269 ( .A(n8127), .B(n5660), .Y(n8171) );
  NOR2X1 U5270 ( .A(n8213), .B(wr_ptr[0]), .Y(n5660) );
  OAI21X1 U5388 ( .A(n5569), .B(n3187), .C(n8254), .Y(n10924) );
  NAND2X1 U5389 ( .A(arr[2622]), .B(n3188), .Y(n8254) );
  OAI21X1 U5391 ( .A(n5571), .B(n3187), .C(n8255), .Y(n10925) );
  NAND2X1 U5392 ( .A(arr[2623]), .B(n3188), .Y(n8255) );
  NAND2X1 U5393 ( .A(n8127), .B(n5703), .Y(n8214) );
  NOR2X1 U5394 ( .A(n8213), .B(n8170), .Y(n5703) );
  NOR2X1 U5396 ( .A(n8084), .B(n7914), .Y(n6215) );
  AND2X1 U5397 ( .A(n7574), .B(wr_ptr[4]), .Y(n7744) );
  OAI21X1 U5400 ( .A(n6896), .B(n8256), .C(n8257), .Y(n10926) );
  NAND2X1 U5401 ( .A(n91), .B(n6895), .Y(n8257) );
  OAI21X1 U5403 ( .A(n6217), .B(n8256), .C(n8258), .Y(n10927) );
  NAND2X1 U5404 ( .A(n90), .B(n6895), .Y(n8258) );
  OAI21X1 U5406 ( .A(n8084), .B(n8256), .C(n8259), .Y(n10928) );
  NAND2X1 U5407 ( .A(n89), .B(n6895), .Y(n8259) );
  OAI21X1 U5409 ( .A(n7914), .B(n8256), .C(n8260), .Y(n10929) );
  NAND2X1 U5410 ( .A(n88), .B(n6895), .Y(n8260) );
  OAI21X1 U5412 ( .A(n8213), .B(n8256), .C(n8261), .Y(n10930) );
  NAND2X1 U5413 ( .A(n87), .B(n6895), .Y(n8261) );
  OAI21X1 U5415 ( .A(n8170), .B(n8256), .C(n8262), .Y(n10931) );
  NAND2X1 U5416 ( .A(n86), .B(n6895), .Y(n8262) );
  NOR2X1 U5417 ( .A(n8263), .B(reset), .Y(n6895) );
  NAND2X1 U5418 ( .A(n8263), .B(n8264), .Y(n8256) );
  OAI21X1 U5421 ( .A(n8266), .B(n8267), .C(n8268), .Y(n10932) );
  AOI22X1 U5422 ( .A(n97), .B(n8269), .C(n2736), .D(n8270), .Y(n8268) );
  OAI21X1 U5424 ( .A(n8266), .B(n8271), .C(n8272), .Y(n10933) );
  AOI22X1 U5425 ( .A(n96), .B(n8269), .C(n2735), .D(n8270), .Y(n8272) );
  OAI21X1 U5426 ( .A(n8266), .B(n8273), .C(n8274), .Y(n10934) );
  AOI22X1 U5427 ( .A(n95), .B(n8269), .C(n2734), .D(n8270), .Y(n8274) );
  OAI21X1 U5428 ( .A(n8266), .B(n8275), .C(n8276), .Y(n10935) );
  AOI22X1 U5429 ( .A(n94), .B(n8269), .C(n2733), .D(n8270), .Y(n8276) );
  OAI21X1 U5430 ( .A(n8266), .B(n8277), .C(n8278), .Y(n10936) );
  AOI22X1 U5431 ( .A(n98), .B(n8269), .C(n2737), .D(n8270), .Y(n8278) );
  OAI21X1 U5433 ( .A(n8266), .B(n8279), .C(n8280), .Y(n10937) );
  AOI22X1 U5434 ( .A(n93), .B(n8269), .C(n2732), .D(n8270), .Y(n8280) );
  OAI21X1 U5435 ( .A(n8266), .B(n8281), .C(n8282), .Y(n10938) );
  AOI22X1 U5436 ( .A(n92), .B(n8269), .C(n2731), .D(n8270), .Y(n8282) );
  NAND3X1 U5438 ( .A(n8266), .B(get), .C(n8284), .Y(n8283) );
  NOR2X1 U5439 ( .A(reset), .B(empty), .Y(n8284) );
  NOR2X1 U5440 ( .A(n8285), .B(n5489), .Y(n8269) );
  OAI21X1 U5442 ( .A(n8265), .B(n5489), .C(n8286), .Y(n8285) );
  NAND3X1 U5443 ( .A(n8287), .B(n8264), .C(n8288), .Y(n8286) );
  NOR2X1 U5444 ( .A(n8289), .B(n8290), .Y(n8288) );
  AOI21X1 U5446 ( .A(n8292), .B(n8293), .C(n8294), .Y(n8291) );
  OAI21X1 U5447 ( .A(empty), .B(n8289), .C(n8264), .Y(n5489) );
  NOR2X1 U5450 ( .A(n8290), .B(full), .Y(n8265) );
  NOR2X1 U5452 ( .A(n8293), .B(n8294), .Y(full) );
  NAND3X1 U5453 ( .A(fillcount[1]), .B(n8281), .C(fillcount[2]), .Y(n8293) );
  NOR2X1 U5454 ( .A(n8294), .B(n8292), .Y(empty) );
  NAND3X1 U5455 ( .A(n8279), .B(n8275), .C(n8281), .Y(n8292) );
  NAND3X1 U5459 ( .A(n8273), .B(n8271), .C(n8295), .Y(n8294) );
  NOR2X1 U5460 ( .A(fillcount[6]), .B(fillcount[5]), .Y(n8295) );
  INVX2 U3 ( .A(n5481), .Y(n8296) );
  INVX2 U5 ( .A(n5484), .Y(n8297) );
  INVX2 U7 ( .A(n5485), .Y(n8298) );
  INVX2 U9 ( .A(n5486), .Y(n8299) );
  INVX2 U11 ( .A(n5487), .Y(n8300) );
  INVX2 U13 ( .A(n5488), .Y(n8301) );
  INVX2 U16 ( .A(n5489), .Y(n5483) );
  INVX2 U5273 ( .A(data_in[0]), .Y(n5491) );
  INVX2 U5276 ( .A(data_in[1]), .Y(n5493) );
  INVX2 U5279 ( .A(data_in[2]), .Y(n5495) );
  INVX2 U5282 ( .A(data_in[3]), .Y(n5497) );
  INVX2 U5285 ( .A(data_in[4]), .Y(n5499) );
  INVX2 U5288 ( .A(data_in[5]), .Y(n5501) );
  INVX2 U5291 ( .A(data_in[6]), .Y(n5503) );
  INVX2 U5294 ( .A(data_in[7]), .Y(n5505) );
  INVX2 U5297 ( .A(data_in[8]), .Y(n5507) );
  INVX2 U5300 ( .A(data_in[9]), .Y(n5509) );
  INVX2 U5303 ( .A(data_in[10]), .Y(n5511) );
  INVX2 U5306 ( .A(data_in[11]), .Y(n5513) );
  INVX2 U5309 ( .A(data_in[12]), .Y(n5515) );
  INVX2 U5312 ( .A(data_in[13]), .Y(n5517) );
  INVX2 U5315 ( .A(data_in[14]), .Y(n5519) );
  INVX2 U5318 ( .A(data_in[15]), .Y(n5521) );
  INVX2 U5321 ( .A(data_in[16]), .Y(n5523) );
  INVX2 U5324 ( .A(data_in[17]), .Y(n5525) );
  INVX2 U5327 ( .A(data_in[18]), .Y(n5527) );
  INVX2 U5330 ( .A(data_in[19]), .Y(n5529) );
  INVX2 U5333 ( .A(data_in[20]), .Y(n5531) );
  INVX2 U5336 ( .A(data_in[21]), .Y(n5533) );
  INVX2 U5339 ( .A(data_in[22]), .Y(n5535) );
  INVX2 U5342 ( .A(data_in[23]), .Y(n5537) );
  INVX2 U5345 ( .A(data_in[24]), .Y(n5539) );
  INVX2 U5348 ( .A(data_in[25]), .Y(n5541) );
  INVX2 U5351 ( .A(data_in[26]), .Y(n5543) );
  INVX2 U5354 ( .A(data_in[27]), .Y(n5545) );
  INVX2 U5357 ( .A(data_in[28]), .Y(n5547) );
  INVX2 U5360 ( .A(data_in[29]), .Y(n5549) );
  INVX2 U5363 ( .A(data_in[30]), .Y(n5551) );
  INVX2 U5366 ( .A(data_in[31]), .Y(n5553) );
  INVX2 U5369 ( .A(data_in[32]), .Y(n5555) );
  INVX2 U5372 ( .A(data_in[33]), .Y(n5557) );
  INVX2 U5375 ( .A(data_in[34]), .Y(n5559) );
  INVX2 U5378 ( .A(data_in[35]), .Y(n5561) );
  INVX2 U5381 ( .A(data_in[36]), .Y(n5563) );
  INVX2 U5384 ( .A(data_in[37]), .Y(n5565) );
  INVX2 U5387 ( .A(data_in[38]), .Y(n5567) );
  INVX2 U5402 ( .A(wr_ptr[5]), .Y(n6896) );
  INVX2 U5405 ( .A(wr_ptr[4]), .Y(n6217) );
  INVX2 U5408 ( .A(wr_ptr[3]), .Y(n8084) );
  INVX2 U5411 ( .A(wr_ptr[2]), .Y(n7914) );
  INVX2 U5414 ( .A(wr_ptr[1]), .Y(n8213) );
  INVX2 U5419 ( .A(n8265), .Y(n8263) );
  INVX2 U5420 ( .A(wr_ptr[0]), .Y(n8170) );
  INVX2 U5437 ( .A(n8283), .Y(n8270) );
  INVX2 U5441 ( .A(n8285), .Y(n8266) );
  INVX2 U5445 ( .A(n8291), .Y(n8287) );
  INVX2 U5448 ( .A(reset), .Y(n8264) );
  INVX2 U5449 ( .A(get), .Y(n8289) );
  INVX2 U5451 ( .A(put), .Y(n8290) );
  INVX2 U5457 ( .A(fillcount[2]), .Y(n8275) );
  INVX2 U5458 ( .A(fillcount[1]), .Y(n8279) );
  INVX2 U5461 ( .A(fillcount[4]), .Y(n8271) );
  INVX2 U5462 ( .A(fillcount[3]), .Y(n8273) );
  FIFO_DEPTH_P26_WIDTH41_DW01_dec_0 sub_55 ( .A(fillcount), .SUM({n2737, n2736, 
        n2735, n2734, n2733, n2732, n2731}) );
  FIFO_DEPTH_P26_WIDTH41_DW01_inc_0 add_54 ( .A({n3555, n17, n16, n15, n14, 
        n13}), .SUM({n2730, n2729, n2728, n2727, n2726, n2725}) );
  FIFO_DEPTH_P26_WIDTH41_DW01_inc_1 add_50 ( .A(fillcount), .SUM({n98, n97, 
        n96, n95, n94, n93, n92}) );
  FIFO_DEPTH_P26_WIDTH41_DW01_inc_2 add_49 ( .A(wr_ptr), .SUM({n91, n90, n89, 
        n88, n87, n86}) );
  BUFX2 U349 ( .A(n5661), .Y(n3533) );
  BUFX2 U682 ( .A(n5661), .Y(n3532) );
  BUFX2 U1015 ( .A(n5661), .Y(n3531) );
  BUFX2 U1348 ( .A(n8042), .Y(n3205) );
  BUFX2 U1682 ( .A(n8214), .Y(n3189) );
  BUFX2 U2015 ( .A(n8042), .Y(n3204) );
  BUFX2 U2348 ( .A(n8214), .Y(n3188) );
  BUFX2 U2681 ( .A(n5661), .Y(n3536) );
  BUFX2 U3016 ( .A(n2923), .Y(n2925) );
  BUFX2 U3349 ( .A(n2923), .Y(n2926) );
  BUFX2 U3682 ( .A(n2922), .Y(n2927) );
  BUFX2 U4015 ( .A(n2922), .Y(n2929) );
  BUFX2 U4349 ( .A(n2922), .Y(n2928) );
  BUFX2 U4683 ( .A(n2921), .Y(n2930) );
  BUFX2 U4685 ( .A(n2921), .Y(n2931) );
  BUFX2 U4686 ( .A(n2920), .Y(n2933) );
  BUFX2 U4687 ( .A(n2921), .Y(n2932) );
  BUFX2 U4688 ( .A(n2920), .Y(n2934) );
  BUFX2 U4689 ( .A(n2920), .Y(n2935) );
  BUFX2 U4690 ( .A(n2919), .Y(n2937) );
  BUFX2 U4691 ( .A(n2919), .Y(n2936) );
  BUFX2 U4692 ( .A(n2919), .Y(n2938) );
  BUFX2 U4693 ( .A(n2918), .Y(n2939) );
  BUFX2 U4694 ( .A(n2918), .Y(n2941) );
  BUFX2 U4695 ( .A(n2918), .Y(n2940) );
  BUFX2 U4696 ( .A(n2917), .Y(n2942) );
  BUFX2 U4697 ( .A(n2917), .Y(n2943) );
  BUFX2 U4698 ( .A(n2916), .Y(n2945) );
  BUFX2 U4699 ( .A(n2917), .Y(n2944) );
  BUFX2 U4700 ( .A(n2916), .Y(n2946) );
  BUFX2 U4701 ( .A(n2916), .Y(n2947) );
  BUFX2 U4702 ( .A(n2915), .Y(n2949) );
  BUFX2 U4703 ( .A(n2915), .Y(n2948) );
  BUFX2 U4704 ( .A(n2915), .Y(n2950) );
  BUFX2 U4705 ( .A(n2914), .Y(n2951) );
  BUFX2 U4706 ( .A(n2914), .Y(n2953) );
  BUFX2 U4707 ( .A(n2914), .Y(n2952) );
  BUFX2 U4708 ( .A(n2913), .Y(n2954) );
  BUFX2 U4709 ( .A(n2913), .Y(n2955) );
  BUFX2 U4710 ( .A(n2912), .Y(n2957) );
  BUFX2 U4711 ( .A(n2913), .Y(n2956) );
  BUFX2 U4712 ( .A(n2912), .Y(n2958) );
  BUFX2 U4713 ( .A(n2912), .Y(n2959) );
  BUFX2 U4714 ( .A(n2911), .Y(n2961) );
  BUFX2 U4715 ( .A(n2911), .Y(n2960) );
  BUFX2 U4716 ( .A(n2911), .Y(n2962) );
  BUFX2 U4717 ( .A(n2910), .Y(n2963) );
  BUFX2 U4718 ( .A(n2910), .Y(n2965) );
  BUFX2 U4719 ( .A(n2910), .Y(n2964) );
  BUFX2 U4720 ( .A(n2909), .Y(n2966) );
  BUFX2 U4721 ( .A(n2909), .Y(n2967) );
  BUFX2 U4722 ( .A(n2908), .Y(n2969) );
  BUFX2 U4723 ( .A(n2909), .Y(n2968) );
  BUFX2 U4724 ( .A(n2908), .Y(n2970) );
  BUFX2 U4725 ( .A(n2908), .Y(n2971) );
  BUFX2 U4726 ( .A(n2907), .Y(n2973) );
  BUFX2 U4727 ( .A(n2907), .Y(n2972) );
  BUFX2 U4728 ( .A(n2907), .Y(n2974) );
  BUFX2 U4729 ( .A(n2906), .Y(n2975) );
  BUFX2 U4730 ( .A(n2906), .Y(n2977) );
  BUFX2 U4731 ( .A(n2906), .Y(n2976) );
  BUFX2 U4732 ( .A(n2905), .Y(n2978) );
  BUFX2 U4733 ( .A(n2905), .Y(n2979) );
  BUFX2 U4734 ( .A(n2904), .Y(n2981) );
  BUFX2 U4735 ( .A(n2905), .Y(n2980) );
  BUFX2 U4736 ( .A(n2904), .Y(n2982) );
  BUFX2 U4737 ( .A(n2904), .Y(n2983) );
  BUFX2 U4738 ( .A(n2903), .Y(n2985) );
  BUFX2 U4739 ( .A(n2903), .Y(n2984) );
  BUFX2 U4740 ( .A(n2903), .Y(n2986) );
  BUFX2 U4741 ( .A(n2902), .Y(n2987) );
  BUFX2 U4742 ( .A(n2902), .Y(n2989) );
  BUFX2 U4743 ( .A(n2902), .Y(n2988) );
  BUFX2 U4744 ( .A(n2901), .Y(n2990) );
  BUFX2 U4745 ( .A(n2901), .Y(n2991) );
  BUFX2 U4746 ( .A(n2900), .Y(n2993) );
  BUFX2 U4747 ( .A(n2901), .Y(n2992) );
  BUFX2 U4748 ( .A(n2900), .Y(n2994) );
  BUFX2 U4749 ( .A(n2900), .Y(n2995) );
  BUFX2 U4750 ( .A(n2899), .Y(n2997) );
  BUFX2 U4751 ( .A(n2899), .Y(n2996) );
  BUFX2 U4752 ( .A(n2899), .Y(n2998) );
  BUFX2 U4753 ( .A(n2898), .Y(n2999) );
  BUFX2 U4754 ( .A(n2898), .Y(n3001) );
  BUFX2 U4755 ( .A(n2898), .Y(n3000) );
  BUFX2 U4756 ( .A(n2897), .Y(n3002) );
  BUFX2 U4757 ( .A(n2897), .Y(n3003) );
  BUFX2 U4758 ( .A(n2896), .Y(n3005) );
  BUFX2 U4759 ( .A(n2897), .Y(n3004) );
  BUFX2 U4760 ( .A(n2896), .Y(n3006) );
  BUFX2 U4761 ( .A(n2896), .Y(n3007) );
  BUFX2 U4762 ( .A(n2895), .Y(n3009) );
  BUFX2 U4768 ( .A(n2895), .Y(n3008) );
  BUFX2 U4769 ( .A(n2895), .Y(n3010) );
  BUFX2 U4770 ( .A(n2894), .Y(n3011) );
  BUFX2 U4771 ( .A(n2894), .Y(n3013) );
  BUFX2 U4772 ( .A(n2894), .Y(n3012) );
  BUFX2 U4773 ( .A(n2893), .Y(n3014) );
  BUFX2 U4774 ( .A(n2893), .Y(n3015) );
  BUFX2 U4775 ( .A(n2892), .Y(n3017) );
  BUFX2 U4776 ( .A(n2893), .Y(n3016) );
  BUFX2 U4777 ( .A(n2892), .Y(n3018) );
  BUFX2 U4778 ( .A(n2892), .Y(n3019) );
  BUFX2 U4779 ( .A(n2891), .Y(n3021) );
  BUFX2 U4780 ( .A(n2891), .Y(n3020) );
  BUFX2 U4781 ( .A(n2891), .Y(n3022) );
  BUFX2 U4782 ( .A(n2890), .Y(n3023) );
  BUFX2 U4783 ( .A(n2890), .Y(n3025) );
  BUFX2 U4784 ( .A(n2890), .Y(n3024) );
  BUFX2 U4785 ( .A(n2889), .Y(n3026) );
  BUFX2 U4786 ( .A(n2889), .Y(n3027) );
  BUFX2 U4787 ( .A(n2888), .Y(n3029) );
  BUFX2 U4788 ( .A(n2889), .Y(n3028) );
  BUFX2 U4789 ( .A(n2888), .Y(n3030) );
  BUFX2 U4790 ( .A(n2888), .Y(n3031) );
  BUFX2 U4791 ( .A(n2923), .Y(n2924) );
  BUFX2 U4792 ( .A(n5575), .Y(n3545) );
  BUFX2 U4793 ( .A(n5575), .Y(n3544) );
  BUFX2 U4794 ( .A(n5575), .Y(n3543) );
  BUFX2 U4795 ( .A(n5618), .Y(n3539) );
  BUFX2 U4796 ( .A(n5618), .Y(n3538) );
  BUFX2 U4797 ( .A(n5618), .Y(n3537) );
  BUFX2 U4798 ( .A(n6940), .Y(n3353) );
  BUFX2 U4799 ( .A(n6940), .Y(n3352) );
  BUFX2 U4800 ( .A(n5490), .Y(n3551) );
  BUFX2 U4801 ( .A(n5490), .Y(n3550) );
  BUFX2 U4802 ( .A(n5490), .Y(n3549) );
  BUFX2 U4803 ( .A(n7915), .Y(n3217) );
  BUFX2 U4804 ( .A(n7958), .Y(n3213) );
  BUFX2 U4805 ( .A(n8000), .Y(n3209) );
  BUFX2 U4806 ( .A(n8085), .Y(n3201) );
  BUFX2 U4807 ( .A(n8128), .Y(n3197) );
  BUFX2 U4808 ( .A(n8171), .Y(n3193) );
  BUFX2 U4809 ( .A(n7915), .Y(n3216) );
  BUFX2 U4810 ( .A(n7958), .Y(n3212) );
  BUFX2 U4811 ( .A(n8000), .Y(n3208) );
  BUFX2 U4812 ( .A(n8085), .Y(n3200) );
  BUFX2 U4813 ( .A(n8128), .Y(n3196) );
  BUFX2 U4814 ( .A(n8171), .Y(n3192) );
  BUFX2 U4815 ( .A(n5490), .Y(n3554) );
  BUFX2 U4816 ( .A(n5575), .Y(n3548) );
  BUFX2 U4817 ( .A(n5618), .Y(n3542) );
  BUFX2 U4818 ( .A(n2887), .Y(n3033) );
  BUFX2 U4819 ( .A(n2887), .Y(n3032) );
  BUFX2 U4820 ( .A(n3110), .Y(n3048) );
  BUFX2 U4821 ( .A(n3110), .Y(n3049) );
  BUFX2 U4822 ( .A(n3110), .Y(n3050) );
  BUFX2 U4823 ( .A(n3111), .Y(n3051) );
  BUFX2 U4824 ( .A(n3111), .Y(n3052) );
  BUFX2 U4825 ( .A(n3111), .Y(n3053) );
  BUFX2 U4826 ( .A(n3112), .Y(n3054) );
  BUFX2 U4827 ( .A(n3112), .Y(n3055) );
  BUFX2 U4828 ( .A(n3112), .Y(n3056) );
  BUFX2 U4829 ( .A(n3113), .Y(n3057) );
  BUFX2 U4830 ( .A(n3113), .Y(n3058) );
  BUFX2 U4831 ( .A(n3113), .Y(n3059) );
  BUFX2 U4832 ( .A(n3114), .Y(n3060) );
  BUFX2 U4833 ( .A(n3114), .Y(n3061) );
  BUFX2 U4834 ( .A(n3114), .Y(n3062) );
  BUFX2 U4835 ( .A(n3115), .Y(n3063) );
  BUFX2 U4836 ( .A(n3115), .Y(n3064) );
  BUFX2 U4837 ( .A(n3115), .Y(n3065) );
  BUFX2 U4838 ( .A(n3116), .Y(n3066) );
  BUFX2 U4839 ( .A(n3116), .Y(n3067) );
  BUFX2 U4840 ( .A(n3116), .Y(n3068) );
  BUFX2 U4841 ( .A(n3117), .Y(n3069) );
  BUFX2 U4842 ( .A(n3117), .Y(n3070) );
  BUFX2 U4843 ( .A(n3117), .Y(n3071) );
  BUFX2 U4844 ( .A(n3118), .Y(n3072) );
  BUFX2 U4845 ( .A(n3118), .Y(n3073) );
  BUFX2 U4851 ( .A(n3118), .Y(n3074) );
  BUFX2 U4852 ( .A(n3119), .Y(n3075) );
  BUFX2 U4853 ( .A(n3119), .Y(n3076) );
  BUFX2 U4854 ( .A(n3119), .Y(n3077) );
  BUFX2 U4855 ( .A(n3120), .Y(n3078) );
  BUFX2 U4856 ( .A(n3120), .Y(n3079) );
  BUFX2 U4857 ( .A(n3120), .Y(n3080) );
  BUFX2 U4858 ( .A(n3121), .Y(n3081) );
  BUFX2 U4859 ( .A(n3121), .Y(n3082) );
  BUFX2 U4860 ( .A(n3121), .Y(n3083) );
  BUFX2 U4861 ( .A(n3122), .Y(n3084) );
  BUFX2 U4862 ( .A(n3122), .Y(n3085) );
  BUFX2 U4863 ( .A(n3122), .Y(n3086) );
  BUFX2 U4864 ( .A(n3123), .Y(n3087) );
  BUFX2 U4865 ( .A(n3123), .Y(n3088) );
  BUFX2 U4866 ( .A(n3123), .Y(n3089) );
  BUFX2 U4867 ( .A(n3124), .Y(n3090) );
  BUFX2 U4868 ( .A(n3124), .Y(n3091) );
  BUFX2 U4869 ( .A(n3124), .Y(n3092) );
  BUFX2 U4870 ( .A(n3125), .Y(n3093) );
  BUFX2 U4871 ( .A(n3125), .Y(n3094) );
  BUFX2 U4872 ( .A(n3125), .Y(n3095) );
  BUFX2 U4873 ( .A(n3126), .Y(n3096) );
  BUFX2 U4874 ( .A(n3126), .Y(n3097) );
  BUFX2 U4875 ( .A(n3126), .Y(n3098) );
  BUFX2 U4876 ( .A(n3157), .Y(n3129) );
  BUFX2 U4877 ( .A(n3157), .Y(n3130) );
  BUFX2 U4878 ( .A(n3157), .Y(n3131) );
  BUFX2 U4879 ( .A(n3158), .Y(n3132) );
  BUFX2 U4880 ( .A(n3158), .Y(n3133) );
  BUFX2 U4881 ( .A(n3158), .Y(n3134) );
  BUFX2 U4882 ( .A(n3159), .Y(n3135) );
  BUFX2 U4883 ( .A(n3159), .Y(n3136) );
  BUFX2 U4884 ( .A(n3159), .Y(n3137) );
  BUFX2 U4885 ( .A(n3160), .Y(n3138) );
  BUFX2 U4886 ( .A(n3160), .Y(n3139) );
  BUFX2 U4887 ( .A(n3160), .Y(n3140) );
  BUFX2 U4888 ( .A(n3161), .Y(n3141) );
  BUFX2 U4889 ( .A(n3161), .Y(n3142) );
  BUFX2 U4890 ( .A(n3161), .Y(n3143) );
  BUFX2 U4891 ( .A(n3162), .Y(n3144) );
  BUFX2 U4892 ( .A(n3162), .Y(n3145) );
  BUFX2 U4893 ( .A(n3162), .Y(n3146) );
  BUFX2 U4894 ( .A(n3163), .Y(n3147) );
  BUFX2 U4895 ( .A(n3163), .Y(n3148) );
  BUFX2 U4896 ( .A(n3163), .Y(n3149) );
  BUFX2 U4897 ( .A(n3164), .Y(n3150) );
  BUFX2 U4898 ( .A(n3164), .Y(n3151) );
  BUFX2 U4899 ( .A(n3164), .Y(n3152) );
  BUFX2 U4900 ( .A(n3165), .Y(n3153) );
  BUFX2 U4901 ( .A(n3165), .Y(n3154) );
  BUFX2 U4902 ( .A(n3165), .Y(n3155) );
  BUFX2 U4903 ( .A(n3046), .Y(n2923) );
  BUFX2 U4904 ( .A(n3046), .Y(n2922) );
  BUFX2 U4905 ( .A(n3046), .Y(n2921) );
  BUFX2 U4906 ( .A(n3045), .Y(n2920) );
  BUFX2 U4907 ( .A(n3045), .Y(n2919) );
  BUFX2 U4908 ( .A(n3045), .Y(n2918) );
  BUFX2 U4909 ( .A(n3044), .Y(n2917) );
  BUFX2 U4910 ( .A(n3044), .Y(n2916) );
  BUFX2 U4911 ( .A(n3044), .Y(n2915) );
  BUFX2 U4912 ( .A(n3043), .Y(n2914) );
  BUFX2 U4913 ( .A(n3043), .Y(n2913) );
  BUFX2 U4914 ( .A(n3043), .Y(n2912) );
  BUFX2 U4915 ( .A(n3042), .Y(n2911) );
  BUFX2 U4916 ( .A(n3042), .Y(n2910) );
  BUFX2 U4917 ( .A(n3042), .Y(n2909) );
  BUFX2 U4918 ( .A(n3041), .Y(n2908) );
  BUFX2 U4919 ( .A(n3041), .Y(n2907) );
  BUFX2 U4920 ( .A(n3041), .Y(n2906) );
  BUFX2 U4921 ( .A(n3040), .Y(n2905) );
  BUFX2 U4922 ( .A(n3040), .Y(n2904) );
  BUFX2 U4923 ( .A(n3040), .Y(n2903) );
  BUFX2 U4924 ( .A(n3039), .Y(n2902) );
  BUFX2 U4925 ( .A(n3039), .Y(n2901) );
  BUFX2 U4926 ( .A(n3039), .Y(n2900) );
  BUFX2 U4927 ( .A(n3038), .Y(n2899) );
  BUFX2 U4928 ( .A(n3038), .Y(n2898) );
  BUFX2 U4934 ( .A(n3038), .Y(n2897) );
  BUFX2 U4935 ( .A(n3037), .Y(n2896) );
  BUFX2 U4936 ( .A(n3037), .Y(n2895) );
  BUFX2 U4937 ( .A(n3037), .Y(n2894) );
  BUFX2 U4938 ( .A(n3036), .Y(n2893) );
  BUFX2 U4939 ( .A(n3036), .Y(n2892) );
  BUFX2 U4940 ( .A(n3036), .Y(n2891) );
  BUFX2 U4941 ( .A(n3035), .Y(n2890) );
  BUFX2 U4942 ( .A(n3035), .Y(n2889) );
  BUFX2 U4943 ( .A(n3035), .Y(n2888) );
  BUFX2 U4944 ( .A(n3127), .Y(n3099) );
  BUFX2 U4945 ( .A(n3127), .Y(n3100) );
  BUFX2 U4946 ( .A(n3127), .Y(n3101) );
  BUFX2 U4947 ( .A(n16), .Y(n3167) );
  BUFX2 U4948 ( .A(n16), .Y(n3168) );
  BUFX2 U4949 ( .A(n16), .Y(n3169) );
  BUFX2 U4950 ( .A(n16), .Y(n3170) );
  BUFX2 U4951 ( .A(n16), .Y(n3171) );
  BUFX2 U4952 ( .A(n16), .Y(n3172) );
  BUFX2 U4953 ( .A(n16), .Y(n3173) );
  BUFX2 U4954 ( .A(n16), .Y(n3174) );
  BUFX2 U4955 ( .A(n16), .Y(n3175) );
  BUFX2 U4956 ( .A(n16), .Y(n3176) );
  BUFX2 U4957 ( .A(n16), .Y(n3177) );
  BUFX2 U4958 ( .A(n16), .Y(n3178) );
  BUFX2 U4959 ( .A(n16), .Y(n3179) );
  BUFX2 U4960 ( .A(n16), .Y(n3166) );
  BUFX2 U4961 ( .A(n3109), .Y(n3047) );
  BUFX2 U4962 ( .A(n3108), .Y(n3109) );
  BUFX2 U4963 ( .A(n3156), .Y(n3128) );
  BUFX2 U4964 ( .A(n15), .Y(n3156) );
  BUFX2 U4965 ( .A(n13), .Y(n3046) );
  BUFX2 U4966 ( .A(n13), .Y(n3045) );
  BUFX2 U4967 ( .A(n13), .Y(n3044) );
  BUFX2 U4968 ( .A(n13), .Y(n3043) );
  BUFX2 U4969 ( .A(n13), .Y(n3042) );
  BUFX2 U4970 ( .A(n13), .Y(n3041) );
  BUFX2 U4971 ( .A(n13), .Y(n3040) );
  BUFX2 U4972 ( .A(n13), .Y(n3039) );
  BUFX2 U4973 ( .A(n13), .Y(n3038) );
  BUFX2 U4974 ( .A(n13), .Y(n3037) );
  BUFX2 U4975 ( .A(n13), .Y(n3036) );
  BUFX2 U4976 ( .A(n13), .Y(n3035) );
  BUFX2 U4977 ( .A(n15), .Y(n3157) );
  BUFX2 U4978 ( .A(n15), .Y(n3158) );
  BUFX2 U4979 ( .A(n15), .Y(n3159) );
  BUFX2 U4980 ( .A(n15), .Y(n3160) );
  BUFX2 U4981 ( .A(n15), .Y(n3161) );
  BUFX2 U4982 ( .A(n15), .Y(n3162) );
  BUFX2 U4983 ( .A(n15), .Y(n3163) );
  BUFX2 U4984 ( .A(n15), .Y(n3164) );
  BUFX2 U4985 ( .A(n15), .Y(n3165) );
  BUFX2 U4986 ( .A(n3108), .Y(n3110) );
  BUFX2 U4987 ( .A(n3108), .Y(n3111) );
  BUFX2 U4988 ( .A(n3107), .Y(n3112) );
  BUFX2 U4989 ( .A(n3107), .Y(n3113) );
  BUFX2 U4990 ( .A(n3107), .Y(n3114) );
  BUFX2 U4991 ( .A(n3106), .Y(n3115) );
  BUFX2 U4992 ( .A(n3106), .Y(n3116) );
  BUFX2 U4993 ( .A(n3106), .Y(n3117) );
  BUFX2 U4994 ( .A(n3105), .Y(n3118) );
  BUFX2 U4995 ( .A(n3105), .Y(n3119) );
  BUFX2 U4996 ( .A(n3105), .Y(n3120) );
  BUFX2 U4997 ( .A(n3104), .Y(n3121) );
  BUFX2 U4998 ( .A(n3104), .Y(n3122) );
  BUFX2 U4999 ( .A(n3104), .Y(n3123) );
  BUFX2 U5000 ( .A(n3103), .Y(n3124) );
  BUFX2 U5001 ( .A(n3103), .Y(n3125) );
  BUFX2 U5002 ( .A(n3103), .Y(n3126) );
  BUFX2 U5003 ( .A(n3034), .Y(n2887) );
  BUFX2 U5004 ( .A(n13), .Y(n3034) );
  INVX2 U5005 ( .A(fillcount[0]), .Y(n8281) );
  AND2X1 U5006 ( .A(arr[2326]), .B(n3218), .Y(n1) );
  AND2X1 U5007 ( .A(arr[2327]), .B(n3218), .Y(n2) );
  AND2X1 U5008 ( .A(arr[2328]), .B(n3218), .Y(n3) );
  AND2X1 U5009 ( .A(arr[2329]), .B(n3218), .Y(n4) );
  AND2X1 U5010 ( .A(arr[2330]), .B(n3218), .Y(n5) );
  AND2X1 U5011 ( .A(arr[2331]), .B(n3218), .Y(n6) );
  AND2X1 U5017 ( .A(arr[2332]), .B(n3218), .Y(n7) );
  AND2X1 U5019 ( .A(arr[2333]), .B(n3218), .Y(n8) );
  AND2X1 U5020 ( .A(arr[2334]), .B(n3218), .Y(n9) );
  AND2X1 U5021 ( .A(arr[2367]), .B(n3214), .Y(n10) );
  AND2X1 U5022 ( .A(arr[2368]), .B(n3214), .Y(n11) );
  AND2X1 U5023 ( .A(arr[2369]), .B(n3214), .Y(n12) );
  AND2X1 U5024 ( .A(arr[2370]), .B(n3214), .Y(n19) );
  AND2X1 U5025 ( .A(arr[2371]), .B(n3214), .Y(n20) );
  AND2X1 U5026 ( .A(arr[2372]), .B(n3214), .Y(n21) );
  AND2X1 U5027 ( .A(arr[2373]), .B(n3214), .Y(n22) );
  AND2X1 U5028 ( .A(arr[2374]), .B(n3214), .Y(n23) );
  AND2X1 U5029 ( .A(arr[2375]), .B(n3214), .Y(n24) );
  AND2X1 U5030 ( .A(arr[2408]), .B(n3210), .Y(n25) );
  AND2X1 U5031 ( .A(arr[2409]), .B(n3210), .Y(n26) );
  AND2X1 U5032 ( .A(arr[2410]), .B(n3210), .Y(n27) );
  AND2X1 U5033 ( .A(arr[2411]), .B(n3210), .Y(n28) );
  AND2X1 U5034 ( .A(arr[2412]), .B(n3210), .Y(n29) );
  AND2X1 U5035 ( .A(arr[2413]), .B(n3210), .Y(n30) );
  AND2X1 U5036 ( .A(arr[2414]), .B(n3210), .Y(n31) );
  AND2X1 U5037 ( .A(arr[2415]), .B(n3210), .Y(n32) );
  AND2X1 U5038 ( .A(arr[2416]), .B(n3210), .Y(n33) );
  AND2X1 U5039 ( .A(arr[2449]), .B(n3206), .Y(n34) );
  AND2X1 U5040 ( .A(arr[2450]), .B(n3206), .Y(n35) );
  AND2X1 U5041 ( .A(arr[2451]), .B(n3206), .Y(n36) );
  AND2X1 U5042 ( .A(arr[2452]), .B(n3206), .Y(n37) );
  AND2X1 U5043 ( .A(arr[2453]), .B(n3206), .Y(n38) );
  AND2X1 U5044 ( .A(arr[2454]), .B(n3206), .Y(n39) );
  AND2X1 U5045 ( .A(arr[2455]), .B(n3206), .Y(n40) );
  AND2X1 U5046 ( .A(arr[2456]), .B(n3206), .Y(n41) );
  AND2X1 U5047 ( .A(arr[2457]), .B(n3206), .Y(n42) );
  AND2X1 U5048 ( .A(arr[2490]), .B(n3202), .Y(n43) );
  AND2X1 U5049 ( .A(arr[2491]), .B(n3202), .Y(n44) );
  AND2X1 U5050 ( .A(arr[2492]), .B(n3202), .Y(n45) );
  AND2X1 U5051 ( .A(arr[2493]), .B(n3202), .Y(n46) );
  AND2X1 U5052 ( .A(arr[2494]), .B(n3202), .Y(n47) );
  AND2X1 U5053 ( .A(arr[2495]), .B(n3202), .Y(n48) );
  AND2X1 U5054 ( .A(arr[2496]), .B(n3202), .Y(n49) );
  AND2X1 U5055 ( .A(arr[2497]), .B(n3202), .Y(n50) );
  AND2X1 U5056 ( .A(arr[2498]), .B(n3202), .Y(n51) );
  AND2X1 U5057 ( .A(arr[2531]), .B(n3198), .Y(n52) );
  AND2X1 U5058 ( .A(arr[2532]), .B(n3198), .Y(n53) );
  AND2X1 U5059 ( .A(arr[2533]), .B(n3198), .Y(n54) );
  AND2X1 U5060 ( .A(arr[2534]), .B(n3198), .Y(n55) );
  AND2X1 U5061 ( .A(arr[2535]), .B(n3198), .Y(n56) );
  AND2X1 U5062 ( .A(arr[2536]), .B(n3198), .Y(n57) );
  AND2X1 U5063 ( .A(arr[2537]), .B(n3198), .Y(n58) );
  AND2X1 U5064 ( .A(arr[2538]), .B(n3198), .Y(n59) );
  AND2X1 U5065 ( .A(arr[2539]), .B(n3198), .Y(n60) );
  AND2X1 U5066 ( .A(arr[2572]), .B(n3194), .Y(n61) );
  AND2X1 U5067 ( .A(arr[2573]), .B(n3194), .Y(n62) );
  AND2X1 U5068 ( .A(arr[2574]), .B(n3194), .Y(n63) );
  AND2X1 U5069 ( .A(arr[2575]), .B(n3194), .Y(n64) );
  AND2X1 U5070 ( .A(arr[2576]), .B(n3194), .Y(n65) );
  AND2X1 U5071 ( .A(arr[2577]), .B(n3194), .Y(n66) );
  AND2X1 U5072 ( .A(arr[2578]), .B(n3194), .Y(n67) );
  AND2X1 U5073 ( .A(arr[2579]), .B(n3194), .Y(n68) );
  AND2X1 U5074 ( .A(arr[2580]), .B(n3194), .Y(n69) );
  AND2X1 U5075 ( .A(arr[2613]), .B(n3190), .Y(n70) );
  AND2X1 U5076 ( .A(arr[2614]), .B(n3190), .Y(n71) );
  AND2X1 U5077 ( .A(arr[2615]), .B(n3190), .Y(n72) );
  AND2X1 U5078 ( .A(arr[2616]), .B(n3190), .Y(n73) );
  AND2X1 U5079 ( .A(arr[2617]), .B(n3190), .Y(n74) );
  AND2X1 U5080 ( .A(arr[2618]), .B(n3190), .Y(n75) );
  AND2X1 U5081 ( .A(arr[2619]), .B(n3190), .Y(n76) );
  AND2X1 U5082 ( .A(arr[2620]), .B(n3190), .Y(n77) );
  AND2X1 U5083 ( .A(arr[2621]), .B(n3190), .Y(n78) );
  AND2X1 U5084 ( .A(arr[2309]), .B(n3217), .Y(n79) );
  AND2X1 U5085 ( .A(arr[2310]), .B(n3217), .Y(n80) );
  AND2X1 U5086 ( .A(arr[2311]), .B(n3217), .Y(n81) );
  AND2X1 U5087 ( .A(arr[2312]), .B(n3217), .Y(n82) );
  AND2X1 U5088 ( .A(arr[2313]), .B(n3217), .Y(n83) );
  AND2X1 U5089 ( .A(arr[2314]), .B(n3217), .Y(n84) );
  AND2X1 U5090 ( .A(arr[2315]), .B(n3217), .Y(n85) );
  AND2X1 U5091 ( .A(arr[2316]), .B(n3217), .Y(n99) );
  AND2X1 U5092 ( .A(arr[2317]), .B(n3217), .Y(n100) );
  AND2X1 U5093 ( .A(arr[2318]), .B(n3217), .Y(n101) );
  AND2X1 U5094 ( .A(arr[2319]), .B(n3217), .Y(n102) );
  AND2X1 U5095 ( .A(arr[2320]), .B(n3217), .Y(n103) );
  AND2X1 U5096 ( .A(arr[2321]), .B(n3217), .Y(n104) );
  AND2X1 U5103 ( .A(arr[2322]), .B(n3217), .Y(n105) );
  AND2X1 U5104 ( .A(arr[2323]), .B(n3217), .Y(n106) );
  AND2X1 U5105 ( .A(arr[2324]), .B(n3217), .Y(n107) );
  AND2X1 U5106 ( .A(arr[2325]), .B(n3217), .Y(n108) );
  AND2X1 U5107 ( .A(arr[2350]), .B(n3213), .Y(n109) );
  AND2X1 U5108 ( .A(arr[2351]), .B(n3213), .Y(n110) );
  AND2X1 U5109 ( .A(arr[2352]), .B(n3213), .Y(n111) );
  AND2X1 U5110 ( .A(arr[2353]), .B(n3213), .Y(n112) );
  AND2X1 U5111 ( .A(arr[2354]), .B(n3213), .Y(n113) );
  AND2X1 U5112 ( .A(arr[2355]), .B(n3213), .Y(n114) );
  AND2X1 U5113 ( .A(arr[2356]), .B(n3213), .Y(n115) );
  AND2X1 U5114 ( .A(arr[2357]), .B(n3213), .Y(n116) );
  AND2X1 U5115 ( .A(arr[2358]), .B(n3213), .Y(n117) );
  AND2X1 U5116 ( .A(arr[2359]), .B(n3213), .Y(n118) );
  AND2X1 U5117 ( .A(arr[2360]), .B(n3213), .Y(n119) );
  AND2X1 U5118 ( .A(arr[2361]), .B(n3213), .Y(n120) );
  AND2X1 U5119 ( .A(arr[2362]), .B(n3213), .Y(n121) );
  AND2X1 U5120 ( .A(arr[2363]), .B(n3213), .Y(n122) );
  AND2X1 U5121 ( .A(arr[2364]), .B(n3213), .Y(n123) );
  AND2X1 U5122 ( .A(arr[2365]), .B(n3213), .Y(n124) );
  AND2X1 U5123 ( .A(arr[2366]), .B(n3213), .Y(n125) );
  AND2X1 U5124 ( .A(arr[2391]), .B(n3209), .Y(n126) );
  AND2X1 U5125 ( .A(arr[2392]), .B(n3209), .Y(n127) );
  AND2X1 U5126 ( .A(arr[2393]), .B(n3209), .Y(n128) );
  AND2X1 U5127 ( .A(arr[2394]), .B(n3209), .Y(n129) );
  AND2X1 U5128 ( .A(arr[2395]), .B(n3209), .Y(n130) );
  AND2X1 U5129 ( .A(arr[2396]), .B(n3209), .Y(n131) );
  AND2X1 U5130 ( .A(arr[2397]), .B(n3209), .Y(n132) );
  AND2X1 U5131 ( .A(arr[2398]), .B(n3209), .Y(n133) );
  AND2X1 U5132 ( .A(arr[2399]), .B(n3209), .Y(n134) );
  AND2X1 U5133 ( .A(arr[2400]), .B(n3209), .Y(n135) );
  AND2X1 U5134 ( .A(arr[2401]), .B(n3209), .Y(n136) );
  AND2X1 U5135 ( .A(arr[2402]), .B(n3209), .Y(n137) );
  AND2X1 U5136 ( .A(arr[2403]), .B(n3209), .Y(n138) );
  AND2X1 U5137 ( .A(arr[2404]), .B(n3209), .Y(n139) );
  AND2X1 U5138 ( .A(arr[2405]), .B(n3209), .Y(n140) );
  AND2X1 U5139 ( .A(arr[2406]), .B(n3209), .Y(n141) );
  AND2X1 U5140 ( .A(arr[2407]), .B(n3209), .Y(n142) );
  AND2X1 U5141 ( .A(arr[2432]), .B(n3205), .Y(n143) );
  AND2X1 U5142 ( .A(arr[2433]), .B(n3205), .Y(n144) );
  AND2X1 U5143 ( .A(arr[2434]), .B(n3205), .Y(n145) );
  AND2X1 U5144 ( .A(arr[2435]), .B(n3205), .Y(n146) );
  AND2X1 U5145 ( .A(arr[2436]), .B(n3205), .Y(n147) );
  AND2X1 U5146 ( .A(arr[2437]), .B(n3205), .Y(n148) );
  AND2X1 U5147 ( .A(arr[2438]), .B(n3205), .Y(n149) );
  AND2X1 U5148 ( .A(arr[2439]), .B(n3205), .Y(n150) );
  AND2X1 U5149 ( .A(arr[2440]), .B(n3205), .Y(n151) );
  AND2X1 U5150 ( .A(arr[2441]), .B(n3205), .Y(n152) );
  AND2X1 U5151 ( .A(arr[2442]), .B(n3205), .Y(n153) );
  AND2X1 U5152 ( .A(arr[2443]), .B(n3205), .Y(n154) );
  AND2X1 U5153 ( .A(arr[2444]), .B(n3205), .Y(n155) );
  AND2X1 U5154 ( .A(arr[2445]), .B(n3205), .Y(n156) );
  AND2X1 U5155 ( .A(arr[2446]), .B(n3205), .Y(n157) );
  AND2X1 U5156 ( .A(arr[2447]), .B(n3205), .Y(n158) );
  AND2X1 U5157 ( .A(arr[2448]), .B(n3205), .Y(n159) );
  AND2X1 U5158 ( .A(arr[2473]), .B(n3201), .Y(n160) );
  AND2X1 U5159 ( .A(arr[2474]), .B(n3201), .Y(n161) );
  AND2X1 U5160 ( .A(arr[2475]), .B(n3201), .Y(n162) );
  AND2X1 U5161 ( .A(arr[2476]), .B(n3201), .Y(n163) );
  AND2X1 U5162 ( .A(arr[2477]), .B(n3201), .Y(n164) );
  AND2X1 U5163 ( .A(arr[2478]), .B(n3201), .Y(n165) );
  AND2X1 U5164 ( .A(arr[2479]), .B(n3201), .Y(n166) );
  AND2X1 U5165 ( .A(arr[2480]), .B(n3201), .Y(n167) );
  AND2X1 U5166 ( .A(arr[2481]), .B(n3201), .Y(n168) );
  AND2X1 U5167 ( .A(arr[2482]), .B(n3201), .Y(n169) );
  AND2X1 U5168 ( .A(arr[2483]), .B(n3201), .Y(n170) );
  AND2X1 U5169 ( .A(arr[2484]), .B(n3201), .Y(n171) );
  AND2X1 U5170 ( .A(arr[2485]), .B(n3201), .Y(n172) );
  AND2X1 U5171 ( .A(arr[2486]), .B(n3201), .Y(n173) );
  AND2X1 U5172 ( .A(arr[2487]), .B(n3201), .Y(n174) );
  AND2X1 U5173 ( .A(arr[2488]), .B(n3201), .Y(n175) );
  AND2X1 U5174 ( .A(arr[2489]), .B(n3201), .Y(n176) );
  AND2X1 U5175 ( .A(arr[2514]), .B(n3197), .Y(n177) );
  AND2X1 U5176 ( .A(arr[2515]), .B(n3197), .Y(n178) );
  AND2X1 U5177 ( .A(arr[2516]), .B(n3197), .Y(n179) );
  AND2X1 U5178 ( .A(arr[2517]), .B(n3197), .Y(n180) );
  AND2X1 U5179 ( .A(arr[2518]), .B(n3197), .Y(n181) );
  AND2X1 U5180 ( .A(arr[2519]), .B(n3197), .Y(n182) );
  AND2X1 U5187 ( .A(arr[2520]), .B(n3197), .Y(n183) );
  AND2X1 U5188 ( .A(arr[2521]), .B(n3197), .Y(n184) );
  AND2X1 U5189 ( .A(arr[2522]), .B(n3197), .Y(n185) );
  AND2X1 U5190 ( .A(arr[2523]), .B(n3197), .Y(n186) );
  AND2X1 U5191 ( .A(arr[2524]), .B(n3197), .Y(n187) );
  AND2X1 U5192 ( .A(arr[2525]), .B(n3197), .Y(n188) );
  AND2X1 U5193 ( .A(arr[2526]), .B(n3197), .Y(n189) );
  AND2X1 U5194 ( .A(arr[2527]), .B(n3197), .Y(n190) );
  AND2X1 U5195 ( .A(arr[2528]), .B(n3197), .Y(n191) );
  AND2X1 U5196 ( .A(arr[2529]), .B(n3197), .Y(n192) );
  AND2X1 U5197 ( .A(arr[2530]), .B(n3197), .Y(n193) );
  AND2X1 U5198 ( .A(arr[2555]), .B(n3193), .Y(n194) );
  AND2X1 U5199 ( .A(arr[2556]), .B(n3193), .Y(n195) );
  AND2X1 U5200 ( .A(arr[2557]), .B(n3193), .Y(n196) );
  AND2X1 U5201 ( .A(arr[2558]), .B(n3193), .Y(n197) );
  AND2X1 U5202 ( .A(arr[2559]), .B(n3193), .Y(n198) );
  AND2X1 U5203 ( .A(arr[2560]), .B(n3193), .Y(n199) );
  AND2X1 U5204 ( .A(arr[2561]), .B(n3193), .Y(n200) );
  AND2X1 U5205 ( .A(arr[2562]), .B(n3193), .Y(n201) );
  AND2X1 U5206 ( .A(arr[2563]), .B(n3193), .Y(n202) );
  AND2X1 U5207 ( .A(arr[2564]), .B(n3193), .Y(n203) );
  AND2X1 U5208 ( .A(arr[2565]), .B(n3193), .Y(n204) );
  AND2X1 U5209 ( .A(arr[2566]), .B(n3193), .Y(n205) );
  AND2X1 U5210 ( .A(arr[2567]), .B(n3193), .Y(n206) );
  AND2X1 U5211 ( .A(arr[2568]), .B(n3193), .Y(n207) );
  AND2X1 U5212 ( .A(arr[2569]), .B(n3193), .Y(n208) );
  AND2X1 U5213 ( .A(arr[2570]), .B(n3193), .Y(n209) );
  AND2X1 U5214 ( .A(arr[2571]), .B(n3193), .Y(n210) );
  AND2X1 U5215 ( .A(arr[2596]), .B(n3189), .Y(n211) );
  AND2X1 U5216 ( .A(arr[2597]), .B(n3189), .Y(n212) );
  AND2X1 U5217 ( .A(arr[2598]), .B(n3189), .Y(n213) );
  AND2X1 U5218 ( .A(arr[2599]), .B(n3189), .Y(n214) );
  AND2X1 U5219 ( .A(arr[2600]), .B(n3189), .Y(n215) );
  AND2X1 U5220 ( .A(arr[2601]), .B(n3189), .Y(n216) );
  AND2X1 U5221 ( .A(arr[2602]), .B(n3189), .Y(n217) );
  AND2X1 U5222 ( .A(arr[2603]), .B(n3189), .Y(n218) );
  AND2X1 U5223 ( .A(arr[2604]), .B(n3189), .Y(n219) );
  AND2X1 U5224 ( .A(arr[2605]), .B(n3189), .Y(n220) );
  AND2X1 U5225 ( .A(arr[2606]), .B(n3189), .Y(n221) );
  AND2X1 U5226 ( .A(arr[2607]), .B(n3189), .Y(n222) );
  AND2X1 U5227 ( .A(arr[2608]), .B(n3189), .Y(n223) );
  AND2X1 U5228 ( .A(arr[2609]), .B(n3189), .Y(n224) );
  AND2X1 U5229 ( .A(arr[2610]), .B(n3189), .Y(n225) );
  AND2X1 U5230 ( .A(arr[2611]), .B(n3189), .Y(n226) );
  AND2X1 U5231 ( .A(arr[2612]), .B(n3189), .Y(n227) );
  AND2X1 U5232 ( .A(arr[2296]), .B(n3216), .Y(n228) );
  AND2X1 U5233 ( .A(arr[2297]), .B(n3216), .Y(n229) );
  AND2X1 U5234 ( .A(arr[2298]), .B(n3216), .Y(n230) );
  AND2X1 U5235 ( .A(arr[2299]), .B(n3216), .Y(n231) );
  AND2X1 U5236 ( .A(arr[2300]), .B(n3216), .Y(n232) );
  AND2X1 U5237 ( .A(arr[2301]), .B(n3216), .Y(n233) );
  AND2X1 U5238 ( .A(arr[2302]), .B(n3216), .Y(n234) );
  AND2X1 U5239 ( .A(arr[2303]), .B(n3216), .Y(n235) );
  AND2X1 U5240 ( .A(arr[2304]), .B(n3216), .Y(n236) );
  AND2X1 U5241 ( .A(arr[2305]), .B(n3216), .Y(n237) );
  AND2X1 U5242 ( .A(arr[2306]), .B(n3216), .Y(n238) );
  AND2X1 U5243 ( .A(arr[2307]), .B(n3216), .Y(n239) );
  AND2X1 U5244 ( .A(arr[2308]), .B(n3216), .Y(n240) );
  AND2X1 U5245 ( .A(arr[2337]), .B(n3212), .Y(n241) );
  AND2X1 U5246 ( .A(arr[2338]), .B(n3212), .Y(n242) );
  AND2X1 U5247 ( .A(arr[2339]), .B(n3212), .Y(n243) );
  AND2X1 U5248 ( .A(arr[2340]), .B(n3212), .Y(n244) );
  AND2X1 U5249 ( .A(arr[2341]), .B(n3212), .Y(n245) );
  AND2X1 U5250 ( .A(arr[2342]), .B(n3212), .Y(n246) );
  AND2X1 U5251 ( .A(arr[2343]), .B(n3212), .Y(n247) );
  AND2X1 U5252 ( .A(arr[2344]), .B(n3212), .Y(n248) );
  AND2X1 U5253 ( .A(arr[2345]), .B(n3212), .Y(n249) );
  AND2X1 U5254 ( .A(arr[2346]), .B(n3212), .Y(n250) );
  AND2X1 U5255 ( .A(arr[2347]), .B(n3212), .Y(n251) );
  AND2X1 U5256 ( .A(arr[2348]), .B(n3212), .Y(n252) );
  AND2X1 U5257 ( .A(arr[2349]), .B(n3212), .Y(n253) );
  AND2X1 U5258 ( .A(arr[2378]), .B(n3208), .Y(n254) );
  AND2X1 U5259 ( .A(arr[2379]), .B(n3208), .Y(n255) );
  AND2X1 U5260 ( .A(arr[2380]), .B(n3208), .Y(n256) );
  AND2X1 U5261 ( .A(arr[2381]), .B(n3208), .Y(n257) );
  AND2X1 U5262 ( .A(arr[2382]), .B(n3208), .Y(n258) );
  AND2X1 U5263 ( .A(arr[2383]), .B(n3208), .Y(n259) );
  AND2X1 U5264 ( .A(arr[2384]), .B(n3208), .Y(n260) );
  AND2X1 U5271 ( .A(arr[2385]), .B(n3208), .Y(n261) );
  AND2X1 U5272 ( .A(arr[2386]), .B(n3208), .Y(n262) );
  AND2X1 U5274 ( .A(arr[2387]), .B(n3208), .Y(n263) );
  AND2X1 U5275 ( .A(arr[2388]), .B(n3208), .Y(n264) );
  AND2X1 U5277 ( .A(arr[2389]), .B(n3208), .Y(n265) );
  AND2X1 U5278 ( .A(arr[2390]), .B(n3208), .Y(n266) );
  AND2X1 U5280 ( .A(arr[2419]), .B(n3204), .Y(n267) );
  AND2X1 U5281 ( .A(arr[2420]), .B(n3204), .Y(n268) );
  AND2X1 U5283 ( .A(arr[2421]), .B(n3204), .Y(n269) );
  AND2X1 U5284 ( .A(arr[2422]), .B(n3204), .Y(n270) );
  AND2X1 U5286 ( .A(arr[2423]), .B(n3204), .Y(n271) );
  AND2X1 U5287 ( .A(arr[2424]), .B(n3204), .Y(n272) );
  AND2X1 U5289 ( .A(arr[2425]), .B(n3204), .Y(n273) );
  AND2X1 U5290 ( .A(arr[2426]), .B(n3204), .Y(n274) );
  AND2X1 U5292 ( .A(arr[2427]), .B(n3204), .Y(n275) );
  AND2X1 U5293 ( .A(arr[2428]), .B(n3204), .Y(n276) );
  AND2X1 U5295 ( .A(arr[2429]), .B(n3204), .Y(n277) );
  AND2X1 U5296 ( .A(arr[2430]), .B(n3204), .Y(n278) );
  AND2X1 U5298 ( .A(arr[2431]), .B(n3204), .Y(n279) );
  AND2X1 U5299 ( .A(arr[2460]), .B(n3200), .Y(n280) );
  AND2X1 U5301 ( .A(arr[2461]), .B(n3200), .Y(n281) );
  AND2X1 U5302 ( .A(arr[2462]), .B(n3200), .Y(n282) );
  AND2X1 U5304 ( .A(arr[2463]), .B(n3200), .Y(n283) );
  AND2X1 U5305 ( .A(arr[2464]), .B(n3200), .Y(n284) );
  AND2X1 U5307 ( .A(arr[2465]), .B(n3200), .Y(n285) );
  AND2X1 U5308 ( .A(arr[2466]), .B(n3200), .Y(n286) );
  AND2X1 U5310 ( .A(arr[2467]), .B(n3200), .Y(n287) );
  AND2X1 U5311 ( .A(arr[2468]), .B(n3200), .Y(n288) );
  AND2X1 U5313 ( .A(arr[2469]), .B(n3200), .Y(n289) );
  AND2X1 U5314 ( .A(arr[2470]), .B(n3200), .Y(n290) );
  AND2X1 U5316 ( .A(arr[2471]), .B(n3200), .Y(n291) );
  AND2X1 U5317 ( .A(arr[2472]), .B(n3200), .Y(n292) );
  AND2X1 U5319 ( .A(arr[2501]), .B(n3196), .Y(n293) );
  AND2X1 U5320 ( .A(arr[2502]), .B(n3196), .Y(n294) );
  AND2X1 U5322 ( .A(arr[2503]), .B(n3196), .Y(n295) );
  AND2X1 U5323 ( .A(arr[2504]), .B(n3196), .Y(n296) );
  AND2X1 U5325 ( .A(arr[2505]), .B(n3196), .Y(n297) );
  AND2X1 U5326 ( .A(arr[2506]), .B(n3196), .Y(n298) );
  AND2X1 U5328 ( .A(arr[2507]), .B(n3196), .Y(n299) );
  AND2X1 U5329 ( .A(arr[2508]), .B(n3196), .Y(n300) );
  AND2X1 U5331 ( .A(arr[2509]), .B(n3196), .Y(n301) );
  AND2X1 U5332 ( .A(arr[2510]), .B(n3196), .Y(n302) );
  AND2X1 U5334 ( .A(arr[2511]), .B(n3196), .Y(n303) );
  AND2X1 U5335 ( .A(arr[2512]), .B(n3196), .Y(n304) );
  AND2X1 U5337 ( .A(arr[2513]), .B(n3196), .Y(n305) );
  AND2X1 U5338 ( .A(arr[2542]), .B(n3192), .Y(n306) );
  AND2X1 U5340 ( .A(arr[2543]), .B(n3192), .Y(n307) );
  AND2X1 U5341 ( .A(arr[2544]), .B(n3192), .Y(n308) );
  AND2X1 U5343 ( .A(arr[2545]), .B(n3192), .Y(n309) );
  AND2X1 U5344 ( .A(arr[2546]), .B(n3192), .Y(n310) );
  AND2X1 U5346 ( .A(arr[2547]), .B(n3192), .Y(n311) );
  AND2X1 U5347 ( .A(arr[2548]), .B(n3192), .Y(n312) );
  AND2X1 U5349 ( .A(arr[2549]), .B(n3192), .Y(n313) );
  AND2X1 U5350 ( .A(arr[2550]), .B(n3192), .Y(n314) );
  AND2X1 U5352 ( .A(arr[2551]), .B(n3192), .Y(n315) );
  AND2X1 U5353 ( .A(arr[2552]), .B(n3192), .Y(n316) );
  AND2X1 U5355 ( .A(arr[2553]), .B(n3192), .Y(n317) );
  AND2X1 U5356 ( .A(arr[2554]), .B(n3192), .Y(n318) );
  AND2X1 U5358 ( .A(arr[2583]), .B(n3188), .Y(n319) );
  AND2X1 U5359 ( .A(arr[2584]), .B(n3188), .Y(n320) );
  AND2X1 U5361 ( .A(arr[2585]), .B(n3188), .Y(n321) );
  AND2X1 U5362 ( .A(arr[2586]), .B(n3188), .Y(n322) );
  AND2X1 U5364 ( .A(arr[2587]), .B(n3188), .Y(n323) );
  AND2X1 U5365 ( .A(arr[2588]), .B(n3188), .Y(n324) );
  AND2X1 U5367 ( .A(arr[2589]), .B(n3188), .Y(n325) );
  AND2X1 U5368 ( .A(arr[2590]), .B(n3188), .Y(n326) );
  AND2X1 U5370 ( .A(arr[2591]), .B(n3188), .Y(n327) );
  AND2X1 U5371 ( .A(arr[2592]), .B(n3188), .Y(n328) );
  AND2X1 U5373 ( .A(arr[2593]), .B(n3188), .Y(n329) );
  AND2X1 U5374 ( .A(arr[2594]), .B(n3188), .Y(n330) );
  AND2X1 U5376 ( .A(arr[2595]), .B(n3188), .Y(n331) );
  INVX2 U5377 ( .A(n3556), .Y(n3555) );
  INVX2 U5379 ( .A(n18), .Y(n3556) );
  BUFX2 U5380 ( .A(n17), .Y(n3181) );
  BUFX2 U5382 ( .A(n17), .Y(n3182) );
  BUFX2 U5383 ( .A(n17), .Y(n3183) );
  BUFX2 U5385 ( .A(n17), .Y(n3184) );
  BUFX2 U5386 ( .A(n17), .Y(n3185) );
  BUFX2 U5390 ( .A(n17), .Y(n3186) );
  BUFX2 U5395 ( .A(n17), .Y(n3180) );
  BUFX2 U5398 ( .A(n14), .Y(n3108) );
  BUFX2 U5399 ( .A(n14), .Y(n3107) );
  BUFX2 U5423 ( .A(n14), .Y(n3106) );
  BUFX2 U5432 ( .A(n14), .Y(n3105) );
  BUFX2 U5456 ( .A(n14), .Y(n3104) );
  BUFX2 U5463 ( .A(n14), .Y(n3103) );
  BUFX2 U5464 ( .A(n3102), .Y(n3127) );
  BUFX2 U5465 ( .A(n14), .Y(n3102) );
  MUX2X1 U5466 ( .B(n333), .A(n334), .S(n3047), .Y(n332) );
  MUX2X1 U5467 ( .B(n336), .A(n337), .S(n3047), .Y(n335) );
  MUX2X1 U5468 ( .B(n339), .A(n340), .S(n3047), .Y(n338) );
  MUX2X1 U5469 ( .B(n342), .A(n343), .S(n3047), .Y(n341) );
  MUX2X1 U5470 ( .B(n345), .A(n346), .S(n3166), .Y(n344) );
  MUX2X1 U5471 ( .B(n348), .A(n349), .S(n3047), .Y(n347) );
  MUX2X1 U5472 ( .B(n351), .A(n352), .S(n3047), .Y(n350) );
  MUX2X1 U5473 ( .B(n354), .A(n355), .S(n3047), .Y(n353) );
  MUX2X1 U5474 ( .B(n357), .A(n358), .S(n3047), .Y(n356) );
  MUX2X1 U5475 ( .B(n360), .A(n361), .S(n3166), .Y(n359) );
  MUX2X1 U5476 ( .B(n363), .A(n364), .S(n3048), .Y(n362) );
  MUX2X1 U5477 ( .B(n366), .A(n367), .S(n3048), .Y(n365) );
  MUX2X1 U5478 ( .B(n369), .A(n370), .S(n3048), .Y(n368) );
  MUX2X1 U5479 ( .B(n372), .A(n373), .S(n3048), .Y(n371) );
  MUX2X1 U5480 ( .B(n375), .A(n376), .S(n3166), .Y(n374) );
  MUX2X1 U5481 ( .B(n378), .A(n379), .S(n3048), .Y(n377) );
  MUX2X1 U5482 ( .B(n381), .A(n382), .S(n3048), .Y(n380) );
  MUX2X1 U5483 ( .B(n384), .A(n385), .S(n3048), .Y(n383) );
  MUX2X1 U5484 ( .B(n387), .A(n388), .S(n3048), .Y(n386) );
  MUX2X1 U5485 ( .B(n390), .A(n391), .S(n3166), .Y(n389) );
  MUX2X1 U5486 ( .B(n392), .A(n393), .S(n18), .Y(data_out[0]) );
  MUX2X1 U5487 ( .B(n395), .A(n396), .S(n3048), .Y(n394) );
  MUX2X1 U5488 ( .B(n398), .A(n399), .S(n3048), .Y(n397) );
  MUX2X1 U5489 ( .B(n401), .A(n402), .S(n3048), .Y(n400) );
  MUX2X1 U5490 ( .B(n404), .A(n405), .S(n3048), .Y(n403) );
  MUX2X1 U5491 ( .B(n407), .A(n408), .S(n3166), .Y(n406) );
  MUX2X1 U5492 ( .B(n410), .A(n411), .S(n3049), .Y(n409) );
  MUX2X1 U5493 ( .B(n413), .A(n414), .S(n3049), .Y(n412) );
  MUX2X1 U5494 ( .B(n416), .A(n417), .S(n3049), .Y(n415) );
  MUX2X1 U5495 ( .B(n419), .A(n420), .S(n3049), .Y(n418) );
  MUX2X1 U5496 ( .B(n422), .A(n423), .S(n3166), .Y(n421) );
  MUX2X1 U5497 ( .B(n425), .A(n426), .S(n3049), .Y(n424) );
  MUX2X1 U5498 ( .B(n428), .A(n429), .S(n3049), .Y(n427) );
  MUX2X1 U5499 ( .B(n431), .A(n432), .S(n3049), .Y(n430) );
  MUX2X1 U5500 ( .B(n434), .A(n435), .S(n3049), .Y(n433) );
  MUX2X1 U5501 ( .B(n437), .A(n438), .S(n3166), .Y(n436) );
  MUX2X1 U5502 ( .B(n440), .A(n441), .S(n3049), .Y(n439) );
  MUX2X1 U5503 ( .B(n443), .A(n444), .S(n3049), .Y(n442) );
  MUX2X1 U5504 ( .B(n446), .A(n447), .S(n3049), .Y(n445) );
  MUX2X1 U5505 ( .B(n449), .A(n450), .S(n3049), .Y(n448) );
  MUX2X1 U5506 ( .B(n452), .A(n453), .S(n3166), .Y(n451) );
  MUX2X1 U5507 ( .B(n454), .A(n455), .S(n18), .Y(data_out[1]) );
  MUX2X1 U5508 ( .B(n457), .A(n458), .S(n3050), .Y(n456) );
  MUX2X1 U5509 ( .B(n460), .A(n461), .S(n3050), .Y(n459) );
  MUX2X1 U5510 ( .B(n463), .A(n464), .S(n3050), .Y(n462) );
  MUX2X1 U5511 ( .B(n466), .A(n467), .S(n3050), .Y(n465) );
  MUX2X1 U5512 ( .B(n469), .A(n470), .S(n3167), .Y(n468) );
  MUX2X1 U5513 ( .B(n472), .A(n473), .S(n3050), .Y(n471) );
  MUX2X1 U5514 ( .B(n475), .A(n476), .S(n3050), .Y(n474) );
  MUX2X1 U5515 ( .B(n478), .A(n479), .S(n3050), .Y(n477) );
  MUX2X1 U5516 ( .B(n481), .A(n482), .S(n3050), .Y(n480) );
  MUX2X1 U5517 ( .B(n484), .A(n485), .S(n3167), .Y(n483) );
  MUX2X1 U5518 ( .B(n487), .A(n488), .S(n3050), .Y(n486) );
  MUX2X1 U5519 ( .B(n490), .A(n491), .S(n3050), .Y(n489) );
  MUX2X1 U5520 ( .B(n493), .A(n494), .S(n3050), .Y(n492) );
  MUX2X1 U5521 ( .B(n496), .A(n497), .S(n3050), .Y(n495) );
  MUX2X1 U5522 ( .B(n499), .A(n500), .S(n3167), .Y(n498) );
  MUX2X1 U5523 ( .B(n502), .A(n503), .S(n3051), .Y(n501) );
  MUX2X1 U5524 ( .B(n505), .A(n506), .S(n3051), .Y(n504) );
  MUX2X1 U5525 ( .B(n508), .A(n509), .S(n3051), .Y(n507) );
  MUX2X1 U5526 ( .B(n511), .A(n512), .S(n3051), .Y(n510) );
  MUX2X1 U5527 ( .B(n514), .A(n515), .S(n3167), .Y(n513) );
  MUX2X1 U5528 ( .B(n516), .A(n517), .S(n18), .Y(data_out[2]) );
  MUX2X1 U5529 ( .B(n519), .A(n520), .S(n3051), .Y(n518) );
  MUX2X1 U5530 ( .B(n522), .A(n523), .S(n3051), .Y(n521) );
  MUX2X1 U5531 ( .B(n525), .A(n526), .S(n3051), .Y(n524) );
  MUX2X1 U5532 ( .B(n528), .A(n529), .S(n3051), .Y(n527) );
  MUX2X1 U5533 ( .B(n531), .A(n532), .S(n3167), .Y(n530) );
  MUX2X1 U5534 ( .B(n534), .A(n535), .S(n3051), .Y(n533) );
  MUX2X1 U5535 ( .B(n537), .A(n538), .S(n3051), .Y(n536) );
  MUX2X1 U5536 ( .B(n540), .A(n541), .S(n3051), .Y(n539) );
  MUX2X1 U5537 ( .B(n543), .A(n544), .S(n3051), .Y(n542) );
  MUX2X1 U5538 ( .B(n546), .A(n547), .S(n3167), .Y(n545) );
  MUX2X1 U5539 ( .B(n549), .A(n550), .S(n3052), .Y(n548) );
  MUX2X1 U5540 ( .B(n552), .A(n553), .S(n3052), .Y(n551) );
  MUX2X1 U5541 ( .B(n555), .A(n556), .S(n3052), .Y(n554) );
  MUX2X1 U5542 ( .B(n558), .A(n559), .S(n3052), .Y(n557) );
  MUX2X1 U5543 ( .B(n561), .A(n562), .S(n3167), .Y(n560) );
  MUX2X1 U5544 ( .B(n564), .A(n565), .S(n3052), .Y(n563) );
  MUX2X1 U5545 ( .B(n567), .A(n568), .S(n3052), .Y(n566) );
  MUX2X1 U5546 ( .B(n570), .A(n571), .S(n3052), .Y(n569) );
  MUX2X1 U5547 ( .B(n573), .A(n574), .S(n3052), .Y(n572) );
  MUX2X1 U5548 ( .B(n576), .A(n577), .S(n3167), .Y(n575) );
  MUX2X1 U5549 ( .B(n578), .A(n579), .S(n18), .Y(data_out[3]) );
  MUX2X1 U5550 ( .B(n581), .A(n582), .S(n3052), .Y(n580) );
  MUX2X1 U5551 ( .B(n584), .A(n585), .S(n3052), .Y(n583) );
  MUX2X1 U5552 ( .B(n587), .A(n588), .S(n3052), .Y(n586) );
  MUX2X1 U5553 ( .B(n590), .A(n591), .S(n3052), .Y(n589) );
  MUX2X1 U5554 ( .B(n593), .A(n594), .S(n3167), .Y(n592) );
  MUX2X1 U5555 ( .B(n596), .A(n597), .S(n3053), .Y(n595) );
  MUX2X1 U5556 ( .B(n599), .A(n600), .S(n3053), .Y(n598) );
  MUX2X1 U5557 ( .B(n602), .A(n603), .S(n3053), .Y(n601) );
  MUX2X1 U5558 ( .B(n605), .A(n606), .S(n3053), .Y(n604) );
  MUX2X1 U5559 ( .B(n608), .A(n609), .S(n3167), .Y(n607) );
  MUX2X1 U5560 ( .B(n611), .A(n612), .S(n3053), .Y(n610) );
  MUX2X1 U5561 ( .B(n614), .A(n615), .S(n3053), .Y(n613) );
  MUX2X1 U5562 ( .B(n617), .A(n618), .S(n3053), .Y(n616) );
  MUX2X1 U5563 ( .B(n620), .A(n621), .S(n3053), .Y(n619) );
  MUX2X1 U5564 ( .B(n623), .A(n624), .S(n3167), .Y(n622) );
  MUX2X1 U5565 ( .B(n626), .A(n627), .S(n3053), .Y(n625) );
  MUX2X1 U5566 ( .B(n629), .A(n630), .S(n3053), .Y(n628) );
  MUX2X1 U5567 ( .B(n632), .A(n633), .S(n3053), .Y(n631) );
  MUX2X1 U5568 ( .B(n635), .A(n636), .S(n3053), .Y(n634) );
  MUX2X1 U5569 ( .B(n638), .A(n639), .S(n3167), .Y(n637) );
  MUX2X1 U5570 ( .B(n640), .A(n641), .S(n18), .Y(data_out[4]) );
  MUX2X1 U5571 ( .B(n643), .A(n644), .S(n3054), .Y(n642) );
  MUX2X1 U5572 ( .B(n646), .A(n647), .S(n3054), .Y(n645) );
  MUX2X1 U5573 ( .B(n649), .A(n650), .S(n3054), .Y(n648) );
  MUX2X1 U5574 ( .B(n652), .A(n653), .S(n3054), .Y(n651) );
  MUX2X1 U5575 ( .B(n655), .A(n656), .S(n3168), .Y(n654) );
  MUX2X1 U5576 ( .B(n658), .A(n659), .S(n3054), .Y(n657) );
  MUX2X1 U5577 ( .B(n661), .A(n662), .S(n3054), .Y(n660) );
  MUX2X1 U5578 ( .B(n664), .A(n665), .S(n3054), .Y(n663) );
  MUX2X1 U5579 ( .B(n667), .A(n668), .S(n3054), .Y(n666) );
  MUX2X1 U5580 ( .B(n670), .A(n671), .S(n3168), .Y(n669) );
  MUX2X1 U5581 ( .B(n673), .A(n674), .S(n3054), .Y(n672) );
  MUX2X1 U5582 ( .B(n676), .A(n677), .S(n3054), .Y(n675) );
  MUX2X1 U5583 ( .B(n679), .A(n680), .S(n3054), .Y(n678) );
  MUX2X1 U5584 ( .B(n682), .A(n683), .S(n3054), .Y(n681) );
  MUX2X1 U5585 ( .B(n685), .A(n686), .S(n3168), .Y(n684) );
  MUX2X1 U5586 ( .B(n688), .A(n689), .S(n3055), .Y(n687) );
  MUX2X1 U5587 ( .B(n691), .A(n692), .S(n3055), .Y(n690) );
  MUX2X1 U5588 ( .B(n694), .A(n695), .S(n3055), .Y(n693) );
  MUX2X1 U5589 ( .B(n697), .A(n698), .S(n3055), .Y(n696) );
  MUX2X1 U5590 ( .B(n700), .A(n701), .S(n3168), .Y(n699) );
  MUX2X1 U5591 ( .B(n702), .A(n703), .S(n18), .Y(data_out[5]) );
  MUX2X1 U5592 ( .B(n705), .A(n706), .S(n3055), .Y(n704) );
  MUX2X1 U5593 ( .B(n708), .A(n709), .S(n3055), .Y(n707) );
  MUX2X1 U5594 ( .B(n711), .A(n712), .S(n3055), .Y(n710) );
  MUX2X1 U5595 ( .B(n714), .A(n715), .S(n3055), .Y(n713) );
  MUX2X1 U5596 ( .B(n717), .A(n718), .S(n3168), .Y(n716) );
  MUX2X1 U5597 ( .B(n720), .A(n721), .S(n3055), .Y(n719) );
  MUX2X1 U5598 ( .B(n723), .A(n724), .S(n3055), .Y(n722) );
  MUX2X1 U5599 ( .B(n726), .A(n727), .S(n3055), .Y(n725) );
  MUX2X1 U5600 ( .B(n729), .A(n730), .S(n3055), .Y(n728) );
  MUX2X1 U5601 ( .B(n732), .A(n733), .S(n3168), .Y(n731) );
  MUX2X1 U5602 ( .B(n735), .A(n736), .S(n3056), .Y(n734) );
  MUX2X1 U5603 ( .B(n738), .A(n739), .S(n3056), .Y(n737) );
  MUX2X1 U5604 ( .B(n741), .A(n742), .S(n3056), .Y(n740) );
  MUX2X1 U5605 ( .B(n744), .A(n745), .S(n3056), .Y(n743) );
  MUX2X1 U5606 ( .B(n747), .A(n748), .S(n3168), .Y(n746) );
  MUX2X1 U5607 ( .B(n750), .A(n751), .S(n3056), .Y(n749) );
  MUX2X1 U5608 ( .B(n753), .A(n754), .S(n3056), .Y(n752) );
  MUX2X1 U5609 ( .B(n756), .A(n757), .S(n3056), .Y(n755) );
  MUX2X1 U5610 ( .B(n759), .A(n760), .S(n3056), .Y(n758) );
  MUX2X1 U5611 ( .B(n762), .A(n763), .S(n3168), .Y(n761) );
  MUX2X1 U5612 ( .B(n764), .A(n765), .S(n18), .Y(data_out[6]) );
  MUX2X1 U5613 ( .B(n767), .A(n768), .S(n3056), .Y(n766) );
  MUX2X1 U5614 ( .B(n770), .A(n771), .S(n3056), .Y(n769) );
  MUX2X1 U5615 ( .B(n773), .A(n774), .S(n3056), .Y(n772) );
  MUX2X1 U5616 ( .B(n776), .A(n777), .S(n3056), .Y(n775) );
  MUX2X1 U5617 ( .B(n779), .A(n780), .S(n3168), .Y(n778) );
  MUX2X1 U5618 ( .B(n782), .A(n783), .S(n3057), .Y(n781) );
  MUX2X1 U5619 ( .B(n785), .A(n786), .S(n3057), .Y(n784) );
  MUX2X1 U5620 ( .B(n788), .A(n789), .S(n3057), .Y(n787) );
  MUX2X1 U5621 ( .B(n791), .A(n792), .S(n3057), .Y(n790) );
  MUX2X1 U5622 ( .B(n794), .A(n795), .S(n3168), .Y(n793) );
  MUX2X1 U5623 ( .B(n797), .A(n798), .S(n3057), .Y(n796) );
  MUX2X1 U5624 ( .B(n800), .A(n801), .S(n3057), .Y(n799) );
  MUX2X1 U5625 ( .B(n803), .A(n804), .S(n3057), .Y(n802) );
  MUX2X1 U5626 ( .B(n806), .A(n807), .S(n3057), .Y(n805) );
  MUX2X1 U5627 ( .B(n809), .A(n810), .S(n3168), .Y(n808) );
  MUX2X1 U5628 ( .B(n812), .A(n813), .S(n3057), .Y(n811) );
  MUX2X1 U5629 ( .B(n815), .A(n816), .S(n3057), .Y(n814) );
  MUX2X1 U5630 ( .B(n818), .A(n819), .S(n3057), .Y(n817) );
  MUX2X1 U5631 ( .B(n821), .A(n822), .S(n3057), .Y(n820) );
  MUX2X1 U5632 ( .B(n824), .A(n825), .S(n3168), .Y(n823) );
  MUX2X1 U5633 ( .B(n826), .A(n827), .S(n18), .Y(data_out[7]) );
  MUX2X1 U5634 ( .B(n829), .A(n830), .S(n3058), .Y(n828) );
  MUX2X1 U5635 ( .B(n832), .A(n833), .S(n3058), .Y(n831) );
  MUX2X1 U5636 ( .B(n835), .A(n836), .S(n3058), .Y(n834) );
  MUX2X1 U5637 ( .B(n838), .A(n839), .S(n3058), .Y(n837) );
  MUX2X1 U5638 ( .B(n841), .A(n842), .S(n3169), .Y(n840) );
  MUX2X1 U5639 ( .B(n844), .A(n845), .S(n3058), .Y(n843) );
  MUX2X1 U5640 ( .B(n847), .A(n848), .S(n3058), .Y(n846) );
  MUX2X1 U5641 ( .B(n850), .A(n851), .S(n3058), .Y(n849) );
  MUX2X1 U5642 ( .B(n853), .A(n854), .S(n3058), .Y(n852) );
  MUX2X1 U5643 ( .B(n856), .A(n857), .S(n3169), .Y(n855) );
  MUX2X1 U5644 ( .B(n859), .A(n860), .S(n3058), .Y(n858) );
  MUX2X1 U5645 ( .B(n862), .A(n863), .S(n3058), .Y(n861) );
  MUX2X1 U5646 ( .B(n865), .A(n866), .S(n3058), .Y(n864) );
  MUX2X1 U5647 ( .B(n868), .A(n869), .S(n3058), .Y(n867) );
  MUX2X1 U5648 ( .B(n871), .A(n872), .S(n3169), .Y(n870) );
  MUX2X1 U5649 ( .B(n874), .A(n875), .S(n3059), .Y(n873) );
  MUX2X1 U5650 ( .B(n877), .A(n878), .S(n3059), .Y(n876) );
  MUX2X1 U5651 ( .B(n880), .A(n881), .S(n3059), .Y(n879) );
  MUX2X1 U5652 ( .B(n883), .A(n884), .S(n3059), .Y(n882) );
  MUX2X1 U5653 ( .B(n886), .A(n887), .S(n3169), .Y(n885) );
  MUX2X1 U5654 ( .B(n888), .A(n889), .S(n18), .Y(data_out[8]) );
  MUX2X1 U5655 ( .B(n891), .A(n892), .S(n3059), .Y(n890) );
  MUX2X1 U5656 ( .B(n894), .A(n895), .S(n3059), .Y(n893) );
  MUX2X1 U5657 ( .B(n897), .A(n898), .S(n3059), .Y(n896) );
  MUX2X1 U5658 ( .B(n900), .A(n901), .S(n3059), .Y(n899) );
  MUX2X1 U5659 ( .B(n903), .A(n904), .S(n3169), .Y(n902) );
  MUX2X1 U5660 ( .B(n906), .A(n907), .S(n3059), .Y(n905) );
  MUX2X1 U5661 ( .B(n909), .A(n910), .S(n3059), .Y(n908) );
  MUX2X1 U5662 ( .B(n912), .A(n913), .S(n3059), .Y(n911) );
  MUX2X1 U5663 ( .B(n915), .A(n916), .S(n3059), .Y(n914) );
  MUX2X1 U5664 ( .B(n918), .A(n919), .S(n3169), .Y(n917) );
  MUX2X1 U5665 ( .B(n921), .A(n922), .S(n3060), .Y(n920) );
  MUX2X1 U5666 ( .B(n924), .A(n925), .S(n3060), .Y(n923) );
  MUX2X1 U5667 ( .B(n927), .A(n928), .S(n3060), .Y(n926) );
  MUX2X1 U5668 ( .B(n930), .A(n931), .S(n3060), .Y(n929) );
  MUX2X1 U5669 ( .B(n933), .A(n934), .S(n3169), .Y(n932) );
  MUX2X1 U5670 ( .B(n936), .A(n937), .S(n3060), .Y(n935) );
  MUX2X1 U5671 ( .B(n939), .A(n940), .S(n3060), .Y(n938) );
  MUX2X1 U5672 ( .B(n942), .A(n943), .S(n3060), .Y(n941) );
  MUX2X1 U5673 ( .B(n945), .A(n946), .S(n3060), .Y(n944) );
  MUX2X1 U5674 ( .B(n948), .A(n949), .S(n3169), .Y(n947) );
  MUX2X1 U5675 ( .B(n950), .A(n951), .S(n18), .Y(data_out[9]) );
  MUX2X1 U5676 ( .B(n953), .A(n954), .S(n3060), .Y(n952) );
  MUX2X1 U5677 ( .B(n956), .A(n957), .S(n3060), .Y(n955) );
  MUX2X1 U5678 ( .B(n959), .A(n960), .S(n3060), .Y(n958) );
  MUX2X1 U5679 ( .B(n962), .A(n963), .S(n3060), .Y(n961) );
  MUX2X1 U5680 ( .B(n965), .A(n966), .S(n3169), .Y(n964) );
  MUX2X1 U5681 ( .B(n968), .A(n969), .S(n3061), .Y(n967) );
  MUX2X1 U5682 ( .B(n971), .A(n972), .S(n3061), .Y(n970) );
  MUX2X1 U5683 ( .B(n974), .A(n975), .S(n3061), .Y(n973) );
  MUX2X1 U5684 ( .B(n977), .A(n978), .S(n3061), .Y(n976) );
  MUX2X1 U5685 ( .B(n980), .A(n981), .S(n3169), .Y(n979) );
  MUX2X1 U5686 ( .B(n983), .A(n984), .S(n3061), .Y(n982) );
  MUX2X1 U5687 ( .B(n986), .A(n987), .S(n3061), .Y(n985) );
  MUX2X1 U5688 ( .B(n989), .A(n990), .S(n3061), .Y(n988) );
  MUX2X1 U5689 ( .B(n992), .A(n993), .S(n3061), .Y(n991) );
  MUX2X1 U5690 ( .B(n995), .A(n996), .S(n3169), .Y(n994) );
  MUX2X1 U5691 ( .B(n998), .A(n999), .S(n3061), .Y(n997) );
  MUX2X1 U5692 ( .B(n1001), .A(n1002), .S(n3061), .Y(n1000) );
  MUX2X1 U5693 ( .B(n1004), .A(n1005), .S(n3061), .Y(n1003) );
  MUX2X1 U5694 ( .B(n1007), .A(n1008), .S(n3061), .Y(n1006) );
  MUX2X1 U5695 ( .B(n1010), .A(n1011), .S(n3169), .Y(n1009) );
  MUX2X1 U5696 ( .B(n1012), .A(n1013), .S(n18), .Y(data_out[10]) );
  MUX2X1 U5697 ( .B(n1015), .A(n1016), .S(n3062), .Y(n1014) );
  MUX2X1 U5698 ( .B(n1018), .A(n1019), .S(n3062), .Y(n1017) );
  MUX2X1 U5699 ( .B(n1021), .A(n1022), .S(n3062), .Y(n1020) );
  MUX2X1 U5700 ( .B(n1024), .A(n1025), .S(n3062), .Y(n1023) );
  MUX2X1 U5701 ( .B(n1027), .A(n1028), .S(n3170), .Y(n1026) );
  MUX2X1 U5702 ( .B(n1030), .A(n1031), .S(n3062), .Y(n1029) );
  MUX2X1 U5703 ( .B(n1033), .A(n1034), .S(n3062), .Y(n1032) );
  MUX2X1 U5704 ( .B(n1036), .A(n1037), .S(n3062), .Y(n1035) );
  MUX2X1 U5705 ( .B(n1039), .A(n1040), .S(n3062), .Y(n1038) );
  MUX2X1 U5706 ( .B(n1042), .A(n1043), .S(n3170), .Y(n1041) );
  MUX2X1 U5707 ( .B(n1045), .A(n1046), .S(n3062), .Y(n1044) );
  MUX2X1 U5708 ( .B(n1048), .A(n1049), .S(n3062), .Y(n1047) );
  MUX2X1 U5709 ( .B(n1051), .A(n1052), .S(n3062), .Y(n1050) );
  MUX2X1 U5710 ( .B(n1054), .A(n1055), .S(n3062), .Y(n1053) );
  MUX2X1 U5711 ( .B(n1057), .A(n1058), .S(n3170), .Y(n1056) );
  MUX2X1 U5712 ( .B(n1060), .A(n1061), .S(n3063), .Y(n1059) );
  MUX2X1 U5713 ( .B(n1063), .A(n1064), .S(n3063), .Y(n1062) );
  MUX2X1 U5714 ( .B(n1066), .A(n1067), .S(n3063), .Y(n1065) );
  MUX2X1 U5715 ( .B(n1069), .A(n1070), .S(n3063), .Y(n1068) );
  MUX2X1 U5716 ( .B(n1072), .A(n1073), .S(n3170), .Y(n1071) );
  MUX2X1 U5717 ( .B(n1074), .A(n1075), .S(n18), .Y(data_out[11]) );
  MUX2X1 U5718 ( .B(n1077), .A(n1078), .S(n3063), .Y(n1076) );
  MUX2X1 U5719 ( .B(n1080), .A(n1081), .S(n3063), .Y(n1079) );
  MUX2X1 U5720 ( .B(n1083), .A(n1084), .S(n3063), .Y(n1082) );
  MUX2X1 U5721 ( .B(n1086), .A(n1087), .S(n3063), .Y(n1085) );
  MUX2X1 U5722 ( .B(n1089), .A(n1090), .S(n3170), .Y(n1088) );
  MUX2X1 U5723 ( .B(n1092), .A(n1093), .S(n3063), .Y(n1091) );
  MUX2X1 U5724 ( .B(n1095), .A(n1096), .S(n3063), .Y(n1094) );
  MUX2X1 U5725 ( .B(n1098), .A(n1099), .S(n3063), .Y(n1097) );
  MUX2X1 U5726 ( .B(n1101), .A(n1102), .S(n3063), .Y(n1100) );
  MUX2X1 U5727 ( .B(n1104), .A(n1105), .S(n3170), .Y(n1103) );
  MUX2X1 U5728 ( .B(n1107), .A(n1108), .S(n3064), .Y(n1106) );
  MUX2X1 U5729 ( .B(n1110), .A(n1111), .S(n3064), .Y(n1109) );
  MUX2X1 U5730 ( .B(n1113), .A(n1114), .S(n3064), .Y(n1112) );
  MUX2X1 U5731 ( .B(n1116), .A(n1117), .S(n3064), .Y(n1115) );
  MUX2X1 U5732 ( .B(n1119), .A(n1120), .S(n3170), .Y(n1118) );
  MUX2X1 U5733 ( .B(n1122), .A(n1123), .S(n3064), .Y(n1121) );
  MUX2X1 U5734 ( .B(n1125), .A(n1126), .S(n3064), .Y(n1124) );
  MUX2X1 U5735 ( .B(n1128), .A(n1129), .S(n3064), .Y(n1127) );
  MUX2X1 U5736 ( .B(n1131), .A(n1132), .S(n3064), .Y(n1130) );
  MUX2X1 U5737 ( .B(n1134), .A(n1135), .S(n3170), .Y(n1133) );
  MUX2X1 U5738 ( .B(n1136), .A(n1137), .S(n18), .Y(data_out[12]) );
  MUX2X1 U5739 ( .B(n1139), .A(n1140), .S(n3064), .Y(n1138) );
  MUX2X1 U5740 ( .B(n1142), .A(n1143), .S(n3064), .Y(n1141) );
  MUX2X1 U5741 ( .B(n1145), .A(n1146), .S(n3064), .Y(n1144) );
  MUX2X1 U5742 ( .B(n1148), .A(n1149), .S(n3064), .Y(n1147) );
  MUX2X1 U5743 ( .B(n1151), .A(n1152), .S(n3170), .Y(n1150) );
  MUX2X1 U5744 ( .B(n1154), .A(n1155), .S(n3065), .Y(n1153) );
  MUX2X1 U5745 ( .B(n1157), .A(n1158), .S(n3065), .Y(n1156) );
  MUX2X1 U5746 ( .B(n1160), .A(n1161), .S(n3065), .Y(n1159) );
  MUX2X1 U5747 ( .B(n1163), .A(n1164), .S(n3065), .Y(n1162) );
  MUX2X1 U5748 ( .B(n1166), .A(n1167), .S(n3170), .Y(n1165) );
  MUX2X1 U5749 ( .B(n1169), .A(n1170), .S(n3065), .Y(n1168) );
  MUX2X1 U5750 ( .B(n1172), .A(n1173), .S(n3065), .Y(n1171) );
  MUX2X1 U5751 ( .B(n1175), .A(n1176), .S(n3065), .Y(n1174) );
  MUX2X1 U5752 ( .B(n1178), .A(n1179), .S(n3065), .Y(n1177) );
  MUX2X1 U5753 ( .B(n1181), .A(n1182), .S(n3170), .Y(n1180) );
  MUX2X1 U5754 ( .B(n1184), .A(n1185), .S(n3065), .Y(n1183) );
  MUX2X1 U5755 ( .B(n1187), .A(n1188), .S(n3065), .Y(n1186) );
  MUX2X1 U5756 ( .B(n1190), .A(n1191), .S(n3065), .Y(n1189) );
  MUX2X1 U5757 ( .B(n1193), .A(n1194), .S(n3065), .Y(n1192) );
  MUX2X1 U5758 ( .B(n1196), .A(n1197), .S(n3170), .Y(n1195) );
  MUX2X1 U5759 ( .B(n1198), .A(n1199), .S(n3555), .Y(data_out[13]) );
  MUX2X1 U5760 ( .B(n1201), .A(n1202), .S(n3066), .Y(n1200) );
  MUX2X1 U5761 ( .B(n1204), .A(n1205), .S(n3066), .Y(n1203) );
  MUX2X1 U5762 ( .B(n1207), .A(n1208), .S(n3066), .Y(n1206) );
  MUX2X1 U5763 ( .B(n1210), .A(n1211), .S(n3066), .Y(n1209) );
  MUX2X1 U5764 ( .B(n1213), .A(n1214), .S(n3171), .Y(n1212) );
  MUX2X1 U5765 ( .B(n1216), .A(n1217), .S(n3066), .Y(n1215) );
  MUX2X1 U5766 ( .B(n1219), .A(n1220), .S(n3066), .Y(n1218) );
  MUX2X1 U5767 ( .B(n1222), .A(n1223), .S(n3066), .Y(n1221) );
  MUX2X1 U5768 ( .B(n1225), .A(n1226), .S(n3066), .Y(n1224) );
  MUX2X1 U5769 ( .B(n1228), .A(n1229), .S(n3171), .Y(n1227) );
  MUX2X1 U5770 ( .B(n1231), .A(n1232), .S(n3066), .Y(n1230) );
  MUX2X1 U5771 ( .B(n1234), .A(n1235), .S(n3066), .Y(n1233) );
  MUX2X1 U5772 ( .B(n1237), .A(n1238), .S(n3066), .Y(n1236) );
  MUX2X1 U5773 ( .B(n1240), .A(n1241), .S(n3066), .Y(n1239) );
  MUX2X1 U5774 ( .B(n1243), .A(n1244), .S(n3171), .Y(n1242) );
  MUX2X1 U5775 ( .B(n1246), .A(n1247), .S(n3067), .Y(n1245) );
  MUX2X1 U5776 ( .B(n1249), .A(n1250), .S(n3067), .Y(n1248) );
  MUX2X1 U5777 ( .B(n1252), .A(n1253), .S(n3067), .Y(n1251) );
  MUX2X1 U5778 ( .B(n1255), .A(n1256), .S(n3067), .Y(n1254) );
  MUX2X1 U5779 ( .B(n1258), .A(n1259), .S(n3171), .Y(n1257) );
  MUX2X1 U5780 ( .B(n1260), .A(n1261), .S(n18), .Y(data_out[14]) );
  MUX2X1 U5781 ( .B(n1263), .A(n1264), .S(n3067), .Y(n1262) );
  MUX2X1 U5782 ( .B(n1266), .A(n1267), .S(n3067), .Y(n1265) );
  MUX2X1 U5783 ( .B(n1269), .A(n1270), .S(n3067), .Y(n1268) );
  MUX2X1 U5784 ( .B(n1272), .A(n1273), .S(n3067), .Y(n1271) );
  MUX2X1 U5785 ( .B(n1275), .A(n1276), .S(n3171), .Y(n1274) );
  MUX2X1 U5786 ( .B(n1278), .A(n1279), .S(n3067), .Y(n1277) );
  MUX2X1 U5787 ( .B(n1281), .A(n1282), .S(n3067), .Y(n1280) );
  MUX2X1 U5788 ( .B(n1284), .A(n1285), .S(n3067), .Y(n1283) );
  MUX2X1 U5789 ( .B(n1287), .A(n1288), .S(n3067), .Y(n1286) );
  MUX2X1 U5790 ( .B(n1290), .A(n1291), .S(n3171), .Y(n1289) );
  MUX2X1 U5791 ( .B(n1293), .A(n1294), .S(n3068), .Y(n1292) );
  MUX2X1 U5792 ( .B(n1296), .A(n1297), .S(n3068), .Y(n1295) );
  MUX2X1 U5793 ( .B(n1299), .A(n1300), .S(n3068), .Y(n1298) );
  MUX2X1 U5794 ( .B(n1302), .A(n1303), .S(n3068), .Y(n1301) );
  MUX2X1 U5795 ( .B(n1305), .A(n1306), .S(n3171), .Y(n1304) );
  MUX2X1 U5796 ( .B(n1308), .A(n1309), .S(n3068), .Y(n1307) );
  MUX2X1 U5797 ( .B(n1311), .A(n1312), .S(n3068), .Y(n1310) );
  MUX2X1 U5798 ( .B(n1314), .A(n1315), .S(n3068), .Y(n1313) );
  MUX2X1 U5799 ( .B(n1317), .A(n1318), .S(n3068), .Y(n1316) );
  MUX2X1 U5800 ( .B(n1320), .A(n1321), .S(n3171), .Y(n1319) );
  MUX2X1 U5801 ( .B(n1322), .A(n1323), .S(n18), .Y(data_out[15]) );
  MUX2X1 U5802 ( .B(n1325), .A(n1326), .S(n3068), .Y(n1324) );
  MUX2X1 U5803 ( .B(n1328), .A(n1329), .S(n3068), .Y(n1327) );
  MUX2X1 U5804 ( .B(n1331), .A(n1332), .S(n3068), .Y(n1330) );
  MUX2X1 U5805 ( .B(n1334), .A(n1335), .S(n3068), .Y(n1333) );
  MUX2X1 U5806 ( .B(n1337), .A(n1338), .S(n3171), .Y(n1336) );
  MUX2X1 U5807 ( .B(n1340), .A(n1341), .S(n3069), .Y(n1339) );
  MUX2X1 U5808 ( .B(n1343), .A(n1344), .S(n3069), .Y(n1342) );
  MUX2X1 U5809 ( .B(n1346), .A(n1347), .S(n3069), .Y(n1345) );
  MUX2X1 U5810 ( .B(n1349), .A(n1350), .S(n3069), .Y(n1348) );
  MUX2X1 U5811 ( .B(n1352), .A(n1353), .S(n3171), .Y(n1351) );
  MUX2X1 U5812 ( .B(n1355), .A(n1356), .S(n3069), .Y(n1354) );
  MUX2X1 U5813 ( .B(n1358), .A(n1359), .S(n3069), .Y(n1357) );
  MUX2X1 U5814 ( .B(n1361), .A(n1362), .S(n3069), .Y(n1360) );
  MUX2X1 U5815 ( .B(n1364), .A(n1365), .S(n3069), .Y(n1363) );
  MUX2X1 U5816 ( .B(n1367), .A(n1368), .S(n3171), .Y(n1366) );
  MUX2X1 U5817 ( .B(n1370), .A(n1371), .S(n3069), .Y(n1369) );
  MUX2X1 U5818 ( .B(n1373), .A(n1374), .S(n3069), .Y(n1372) );
  MUX2X1 U5819 ( .B(n1376), .A(n1377), .S(n3069), .Y(n1375) );
  MUX2X1 U5820 ( .B(n1379), .A(n1380), .S(n3069), .Y(n1378) );
  MUX2X1 U5821 ( .B(n1382), .A(n1383), .S(n3171), .Y(n1381) );
  MUX2X1 U5822 ( .B(n1384), .A(n1385), .S(n18), .Y(data_out[16]) );
  MUX2X1 U5823 ( .B(n1387), .A(n1388), .S(n3070), .Y(n1386) );
  MUX2X1 U5824 ( .B(n1390), .A(n1391), .S(n3070), .Y(n1389) );
  MUX2X1 U5825 ( .B(n1393), .A(n1394), .S(n3070), .Y(n1392) );
  MUX2X1 U5826 ( .B(n1396), .A(n1397), .S(n3070), .Y(n1395) );
  MUX2X1 U5827 ( .B(n1399), .A(n1400), .S(n3172), .Y(n1398) );
  MUX2X1 U5828 ( .B(n1402), .A(n1403), .S(n3070), .Y(n1401) );
  MUX2X1 U5829 ( .B(n1405), .A(n1406), .S(n3070), .Y(n1404) );
  MUX2X1 U5830 ( .B(n1408), .A(n1409), .S(n3070), .Y(n1407) );
  MUX2X1 U5831 ( .B(n1411), .A(n1412), .S(n3070), .Y(n1410) );
  MUX2X1 U5832 ( .B(n1414), .A(n1415), .S(n3172), .Y(n1413) );
  MUX2X1 U5833 ( .B(n1417), .A(n1418), .S(n3070), .Y(n1416) );
  MUX2X1 U5834 ( .B(n1420), .A(n1421), .S(n3070), .Y(n1419) );
  MUX2X1 U5835 ( .B(n1423), .A(n1424), .S(n3070), .Y(n1422) );
  MUX2X1 U5836 ( .B(n1426), .A(n1427), .S(n3070), .Y(n1425) );
  MUX2X1 U5837 ( .B(n1429), .A(n1430), .S(n3172), .Y(n1428) );
  MUX2X1 U5838 ( .B(n1432), .A(n1433), .S(n3071), .Y(n1431) );
  MUX2X1 U5839 ( .B(n1435), .A(n1436), .S(n3071), .Y(n1434) );
  MUX2X1 U5840 ( .B(n1438), .A(n1439), .S(n3071), .Y(n1437) );
  MUX2X1 U5841 ( .B(n1441), .A(n1442), .S(n3071), .Y(n1440) );
  MUX2X1 U5842 ( .B(n1444), .A(n1445), .S(n3172), .Y(n1443) );
  MUX2X1 U5843 ( .B(n1446), .A(n1447), .S(n18), .Y(data_out[17]) );
  MUX2X1 U5844 ( .B(n1449), .A(n1450), .S(n3071), .Y(n1448) );
  MUX2X1 U5845 ( .B(n1452), .A(n1453), .S(n3071), .Y(n1451) );
  MUX2X1 U5846 ( .B(n1455), .A(n1456), .S(n3071), .Y(n1454) );
  MUX2X1 U5847 ( .B(n1458), .A(n1459), .S(n3071), .Y(n1457) );
  MUX2X1 U5848 ( .B(n1461), .A(n1462), .S(n3172), .Y(n1460) );
  MUX2X1 U5849 ( .B(n1464), .A(n1465), .S(n3071), .Y(n1463) );
  MUX2X1 U5850 ( .B(n1467), .A(n1468), .S(n3071), .Y(n1466) );
  MUX2X1 U5851 ( .B(n1470), .A(n1471), .S(n3071), .Y(n1469) );
  MUX2X1 U5852 ( .B(n1473), .A(n1474), .S(n3071), .Y(n1472) );
  MUX2X1 U5853 ( .B(n1476), .A(n1477), .S(n3172), .Y(n1475) );
  MUX2X1 U5854 ( .B(n1479), .A(n1480), .S(n3072), .Y(n1478) );
  MUX2X1 U5855 ( .B(n1482), .A(n1483), .S(n3072), .Y(n1481) );
  MUX2X1 U5856 ( .B(n1485), .A(n1486), .S(n3072), .Y(n1484) );
  MUX2X1 U5857 ( .B(n1488), .A(n1489), .S(n3072), .Y(n1487) );
  MUX2X1 U5858 ( .B(n1491), .A(n1492), .S(n3172), .Y(n1490) );
  MUX2X1 U5859 ( .B(n1494), .A(n1495), .S(n3072), .Y(n1493) );
  MUX2X1 U5860 ( .B(n1497), .A(n1498), .S(n3072), .Y(n1496) );
  MUX2X1 U5861 ( .B(n1500), .A(n1501), .S(n3072), .Y(n1499) );
  MUX2X1 U5862 ( .B(n1503), .A(n1504), .S(n3072), .Y(n1502) );
  MUX2X1 U5863 ( .B(n1506), .A(n1507), .S(n3172), .Y(n1505) );
  MUX2X1 U5864 ( .B(n1508), .A(n1509), .S(n18), .Y(data_out[18]) );
  MUX2X1 U5865 ( .B(n1511), .A(n1512), .S(n3072), .Y(n1510) );
  MUX2X1 U5866 ( .B(n1514), .A(n1515), .S(n3072), .Y(n1513) );
  MUX2X1 U5867 ( .B(n1517), .A(n1518), .S(n3072), .Y(n1516) );
  MUX2X1 U5868 ( .B(n1520), .A(n1521), .S(n3072), .Y(n1519) );
  MUX2X1 U5869 ( .B(n1523), .A(n1524), .S(n3172), .Y(n1522) );
  MUX2X1 U5870 ( .B(n1526), .A(n1527), .S(n3073), .Y(n1525) );
  MUX2X1 U5871 ( .B(n1529), .A(n1530), .S(n3073), .Y(n1528) );
  MUX2X1 U5872 ( .B(n1532), .A(n1533), .S(n3073), .Y(n1531) );
  MUX2X1 U5873 ( .B(n1535), .A(n1536), .S(n3073), .Y(n1534) );
  MUX2X1 U5874 ( .B(n1538), .A(n1539), .S(n3172), .Y(n1537) );
  MUX2X1 U5875 ( .B(n1541), .A(n1542), .S(n3073), .Y(n1540) );
  MUX2X1 U5876 ( .B(n1544), .A(n1545), .S(n3073), .Y(n1543) );
  MUX2X1 U5877 ( .B(n1547), .A(n1548), .S(n3073), .Y(n1546) );
  MUX2X1 U5878 ( .B(n1550), .A(n1551), .S(n3073), .Y(n1549) );
  MUX2X1 U5879 ( .B(n1553), .A(n1554), .S(n3172), .Y(n1552) );
  MUX2X1 U5880 ( .B(n1556), .A(n1557), .S(n3073), .Y(n1555) );
  MUX2X1 U5881 ( .B(n1559), .A(n1560), .S(n3073), .Y(n1558) );
  MUX2X1 U5882 ( .B(n1562), .A(n1563), .S(n3073), .Y(n1561) );
  MUX2X1 U5883 ( .B(n1565), .A(n1566), .S(n3073), .Y(n1564) );
  MUX2X1 U5884 ( .B(n1568), .A(n1569), .S(n3172), .Y(n1567) );
  MUX2X1 U5885 ( .B(n1570), .A(n1571), .S(n18), .Y(data_out[19]) );
  MUX2X1 U5886 ( .B(n1573), .A(n1574), .S(n3074), .Y(n1572) );
  MUX2X1 U5887 ( .B(n1576), .A(n1577), .S(n3074), .Y(n1575) );
  MUX2X1 U5888 ( .B(n1579), .A(n1580), .S(n3074), .Y(n1578) );
  MUX2X1 U5889 ( .B(n1582), .A(n1583), .S(n3074), .Y(n1581) );
  MUX2X1 U5890 ( .B(n1585), .A(n1586), .S(n3173), .Y(n1584) );
  MUX2X1 U5891 ( .B(n1588), .A(n1589), .S(n3074), .Y(n1587) );
  MUX2X1 U5892 ( .B(n1591), .A(n1592), .S(n3074), .Y(n1590) );
  MUX2X1 U5893 ( .B(n1594), .A(n1595), .S(n3074), .Y(n1593) );
  MUX2X1 U5894 ( .B(n1597), .A(n1598), .S(n3074), .Y(n1596) );
  MUX2X1 U5895 ( .B(n1600), .A(n1601), .S(n3173), .Y(n1599) );
  MUX2X1 U5896 ( .B(n1603), .A(n1604), .S(n3074), .Y(n1602) );
  MUX2X1 U5897 ( .B(n1606), .A(n1607), .S(n3074), .Y(n1605) );
  MUX2X1 U5898 ( .B(n1609), .A(n1610), .S(n3074), .Y(n1608) );
  MUX2X1 U5899 ( .B(n1612), .A(n1613), .S(n3074), .Y(n1611) );
  MUX2X1 U5900 ( .B(n1615), .A(n1616), .S(n3173), .Y(n1614) );
  MUX2X1 U5901 ( .B(n1618), .A(n1619), .S(n3075), .Y(n1617) );
  MUX2X1 U5902 ( .B(n1621), .A(n1622), .S(n3075), .Y(n1620) );
  MUX2X1 U5903 ( .B(n1624), .A(n1625), .S(n3075), .Y(n1623) );
  MUX2X1 U5904 ( .B(n1627), .A(n1628), .S(n3075), .Y(n1626) );
  MUX2X1 U5905 ( .B(n1630), .A(n1631), .S(n3173), .Y(n1629) );
  MUX2X1 U5906 ( .B(n1632), .A(n1633), .S(n18), .Y(data_out[20]) );
  MUX2X1 U5907 ( .B(n1635), .A(n1636), .S(n3075), .Y(n1634) );
  MUX2X1 U5908 ( .B(n1638), .A(n1639), .S(n3075), .Y(n1637) );
  MUX2X1 U5909 ( .B(n1641), .A(n1642), .S(n3075), .Y(n1640) );
  MUX2X1 U5910 ( .B(n1644), .A(n1645), .S(n3075), .Y(n1643) );
  MUX2X1 U5911 ( .B(n1647), .A(n1648), .S(n3173), .Y(n1646) );
  MUX2X1 U5912 ( .B(n1650), .A(n1651), .S(n3075), .Y(n1649) );
  MUX2X1 U5913 ( .B(n1653), .A(n1654), .S(n3075), .Y(n1652) );
  MUX2X1 U5914 ( .B(n1656), .A(n1657), .S(n3075), .Y(n1655) );
  MUX2X1 U5915 ( .B(n1659), .A(n1660), .S(n3075), .Y(n1658) );
  MUX2X1 U5916 ( .B(n1662), .A(n1663), .S(n3173), .Y(n1661) );
  MUX2X1 U5917 ( .B(n1665), .A(n1666), .S(n3076), .Y(n1664) );
  MUX2X1 U5918 ( .B(n1668), .A(n1669), .S(n3076), .Y(n1667) );
  MUX2X1 U5919 ( .B(n1671), .A(n1672), .S(n3076), .Y(n1670) );
  MUX2X1 U5920 ( .B(n1674), .A(n1675), .S(n3076), .Y(n1673) );
  MUX2X1 U5921 ( .B(n1677), .A(n1678), .S(n3173), .Y(n1676) );
  MUX2X1 U5922 ( .B(n1680), .A(n1681), .S(n3076), .Y(n1679) );
  MUX2X1 U5923 ( .B(n1683), .A(n1684), .S(n3076), .Y(n1682) );
  MUX2X1 U5924 ( .B(n1686), .A(n1687), .S(n3076), .Y(n1685) );
  MUX2X1 U5925 ( .B(n1689), .A(n1690), .S(n3076), .Y(n1688) );
  MUX2X1 U5926 ( .B(n1692), .A(n1693), .S(n3173), .Y(n1691) );
  MUX2X1 U5927 ( .B(n1694), .A(n1695), .S(n18), .Y(data_out[21]) );
  MUX2X1 U5928 ( .B(n1697), .A(n1698), .S(n3076), .Y(n1696) );
  MUX2X1 U5929 ( .B(n1700), .A(n1701), .S(n3076), .Y(n1699) );
  MUX2X1 U5930 ( .B(n1703), .A(n1704), .S(n3076), .Y(n1702) );
  MUX2X1 U5931 ( .B(n1706), .A(n1707), .S(n3076), .Y(n1705) );
  MUX2X1 U5932 ( .B(n1709), .A(n1710), .S(n3173), .Y(n1708) );
  MUX2X1 U5933 ( .B(n1712), .A(n1713), .S(n3077), .Y(n1711) );
  MUX2X1 U5934 ( .B(n1715), .A(n1716), .S(n3077), .Y(n1714) );
  MUX2X1 U5935 ( .B(n1718), .A(n1719), .S(n3077), .Y(n1717) );
  MUX2X1 U5936 ( .B(n1721), .A(n1722), .S(n3077), .Y(n1720) );
  MUX2X1 U5937 ( .B(n1724), .A(n1725), .S(n3173), .Y(n1723) );
  MUX2X1 U5938 ( .B(n1727), .A(n1728), .S(n3077), .Y(n1726) );
  MUX2X1 U5939 ( .B(n1730), .A(n1731), .S(n3077), .Y(n1729) );
  MUX2X1 U5940 ( .B(n1733), .A(n1734), .S(n3077), .Y(n1732) );
  MUX2X1 U5941 ( .B(n1736), .A(n1737), .S(n3077), .Y(n1735) );
  MUX2X1 U5942 ( .B(n1739), .A(n1740), .S(n3173), .Y(n1738) );
  MUX2X1 U5943 ( .B(n1742), .A(n1743), .S(n3077), .Y(n1741) );
  MUX2X1 U5944 ( .B(n1745), .A(n1746), .S(n3077), .Y(n1744) );
  MUX2X1 U5945 ( .B(n1748), .A(n1749), .S(n3077), .Y(n1747) );
  MUX2X1 U5946 ( .B(n1751), .A(n1752), .S(n3077), .Y(n1750) );
  MUX2X1 U5947 ( .B(n1754), .A(n1755), .S(n3173), .Y(n1753) );
  MUX2X1 U5948 ( .B(n1756), .A(n1757), .S(n18), .Y(data_out[22]) );
  MUX2X1 U5949 ( .B(n1759), .A(n1760), .S(n3078), .Y(n1758) );
  MUX2X1 U5950 ( .B(n1762), .A(n1763), .S(n3078), .Y(n1761) );
  MUX2X1 U5951 ( .B(n1765), .A(n1766), .S(n3078), .Y(n1764) );
  MUX2X1 U5952 ( .B(n1768), .A(n1769), .S(n3078), .Y(n1767) );
  MUX2X1 U5953 ( .B(n1771), .A(n1772), .S(n3174), .Y(n1770) );
  MUX2X1 U5954 ( .B(n1774), .A(n1775), .S(n3078), .Y(n1773) );
  MUX2X1 U5955 ( .B(n1777), .A(n1778), .S(n3078), .Y(n1776) );
  MUX2X1 U5956 ( .B(n1780), .A(n1781), .S(n3078), .Y(n1779) );
  MUX2X1 U5957 ( .B(n1783), .A(n1784), .S(n3078), .Y(n1782) );
  MUX2X1 U5958 ( .B(n1786), .A(n1787), .S(n3174), .Y(n1785) );
  MUX2X1 U5959 ( .B(n1789), .A(n1790), .S(n3078), .Y(n1788) );
  MUX2X1 U5960 ( .B(n1792), .A(n1793), .S(n3078), .Y(n1791) );
  MUX2X1 U5961 ( .B(n1795), .A(n1796), .S(n3078), .Y(n1794) );
  MUX2X1 U5962 ( .B(n1798), .A(n1799), .S(n3078), .Y(n1797) );
  MUX2X1 U5963 ( .B(n1801), .A(n1802), .S(n3174), .Y(n1800) );
  MUX2X1 U5964 ( .B(n1804), .A(n1805), .S(n3079), .Y(n1803) );
  MUX2X1 U5965 ( .B(n1807), .A(n1808), .S(n3079), .Y(n1806) );
  MUX2X1 U5966 ( .B(n1810), .A(n1811), .S(n3079), .Y(n1809) );
  MUX2X1 U5967 ( .B(n1813), .A(n1814), .S(n3079), .Y(n1812) );
  MUX2X1 U5968 ( .B(n1816), .A(n1817), .S(n3174), .Y(n1815) );
  MUX2X1 U5969 ( .B(n1818), .A(n1819), .S(n18), .Y(data_out[23]) );
  MUX2X1 U5970 ( .B(n1821), .A(n1822), .S(n3079), .Y(n1820) );
  MUX2X1 U5971 ( .B(n1824), .A(n1825), .S(n3079), .Y(n1823) );
  MUX2X1 U5972 ( .B(n1827), .A(n1828), .S(n3079), .Y(n1826) );
  MUX2X1 U5973 ( .B(n1830), .A(n1831), .S(n3079), .Y(n1829) );
  MUX2X1 U5974 ( .B(n1833), .A(n1834), .S(n3174), .Y(n1832) );
  MUX2X1 U5975 ( .B(n1836), .A(n1837), .S(n3079), .Y(n1835) );
  MUX2X1 U5976 ( .B(n1839), .A(n1840), .S(n3079), .Y(n1838) );
  MUX2X1 U5977 ( .B(n1842), .A(n1843), .S(n3079), .Y(n1841) );
  MUX2X1 U5978 ( .B(n1845), .A(n1846), .S(n3079), .Y(n1844) );
  MUX2X1 U5979 ( .B(n1848), .A(n1849), .S(n3174), .Y(n1847) );
  MUX2X1 U5980 ( .B(n1851), .A(n1852), .S(n3080), .Y(n1850) );
  MUX2X1 U5981 ( .B(n1854), .A(n1855), .S(n3080), .Y(n1853) );
  MUX2X1 U5982 ( .B(n1857), .A(n1858), .S(n3080), .Y(n1856) );
  MUX2X1 U5983 ( .B(n1860), .A(n1861), .S(n3080), .Y(n1859) );
  MUX2X1 U5984 ( .B(n1863), .A(n1864), .S(n3174), .Y(n1862) );
  MUX2X1 U5985 ( .B(n1866), .A(n1867), .S(n3080), .Y(n1865) );
  MUX2X1 U5986 ( .B(n1869), .A(n1870), .S(n3080), .Y(n1868) );
  MUX2X1 U5987 ( .B(n1872), .A(n1873), .S(n3080), .Y(n1871) );
  MUX2X1 U5988 ( .B(n1875), .A(n1876), .S(n3080), .Y(n1874) );
  MUX2X1 U5989 ( .B(n1878), .A(n1879), .S(n3174), .Y(n1877) );
  MUX2X1 U5990 ( .B(n1880), .A(n1881), .S(n18), .Y(data_out[24]) );
  MUX2X1 U5991 ( .B(n1883), .A(n1884), .S(n3080), .Y(n1882) );
  MUX2X1 U5992 ( .B(n1886), .A(n1887), .S(n3080), .Y(n1885) );
  MUX2X1 U5993 ( .B(n1889), .A(n1890), .S(n3080), .Y(n1888) );
  MUX2X1 U5994 ( .B(n1892), .A(n1893), .S(n3080), .Y(n1891) );
  MUX2X1 U5995 ( .B(n1895), .A(n1896), .S(n3174), .Y(n1894) );
  MUX2X1 U5996 ( .B(n1898), .A(n1899), .S(n3081), .Y(n1897) );
  MUX2X1 U5997 ( .B(n1901), .A(n1902), .S(n3081), .Y(n1900) );
  MUX2X1 U5998 ( .B(n1904), .A(n1905), .S(n3081), .Y(n1903) );
  MUX2X1 U5999 ( .B(n1907), .A(n1908), .S(n3081), .Y(n1906) );
  MUX2X1 U6000 ( .B(n1910), .A(n1911), .S(n3174), .Y(n1909) );
  MUX2X1 U6001 ( .B(n1913), .A(n1914), .S(n3081), .Y(n1912) );
  MUX2X1 U6002 ( .B(n1916), .A(n1917), .S(n3081), .Y(n1915) );
  MUX2X1 U6003 ( .B(n1919), .A(n1920), .S(n3081), .Y(n1918) );
  MUX2X1 U6004 ( .B(n1922), .A(n1923), .S(n3081), .Y(n1921) );
  MUX2X1 U6005 ( .B(n1925), .A(n1926), .S(n3174), .Y(n1924) );
  MUX2X1 U6006 ( .B(n1928), .A(n1929), .S(n3081), .Y(n1927) );
  MUX2X1 U6007 ( .B(n1931), .A(n1932), .S(n3081), .Y(n1930) );
  MUX2X1 U6008 ( .B(n1934), .A(n1935), .S(n3081), .Y(n1933) );
  MUX2X1 U6009 ( .B(n1937), .A(n1938), .S(n3081), .Y(n1936) );
  MUX2X1 U6010 ( .B(n1940), .A(n1941), .S(n3174), .Y(n1939) );
  MUX2X1 U6011 ( .B(n1942), .A(n1943), .S(n18), .Y(data_out[25]) );
  MUX2X1 U6012 ( .B(n1945), .A(n1946), .S(n3082), .Y(n1944) );
  MUX2X1 U6013 ( .B(n1948), .A(n1949), .S(n3082), .Y(n1947) );
  MUX2X1 U6014 ( .B(n1951), .A(n1952), .S(n3082), .Y(n1950) );
  MUX2X1 U6015 ( .B(n1954), .A(n1955), .S(n3082), .Y(n1953) );
  MUX2X1 U6016 ( .B(n1957), .A(n1958), .S(n3175), .Y(n1956) );
  MUX2X1 U6017 ( .B(n1960), .A(n1961), .S(n3082), .Y(n1959) );
  MUX2X1 U6018 ( .B(n1963), .A(n1964), .S(n3082), .Y(n1962) );
  MUX2X1 U6019 ( .B(n1966), .A(n1967), .S(n3082), .Y(n1965) );
  MUX2X1 U6020 ( .B(n1969), .A(n1970), .S(n3082), .Y(n1968) );
  MUX2X1 U6021 ( .B(n1972), .A(n1973), .S(n3175), .Y(n1971) );
  MUX2X1 U6022 ( .B(n1975), .A(n1976), .S(n3082), .Y(n1974) );
  MUX2X1 U6023 ( .B(n1978), .A(n1979), .S(n3082), .Y(n1977) );
  MUX2X1 U6024 ( .B(n1981), .A(n1982), .S(n3082), .Y(n1980) );
  MUX2X1 U6025 ( .B(n1984), .A(n1985), .S(n3082), .Y(n1983) );
  MUX2X1 U6026 ( .B(n1987), .A(n1988), .S(n3175), .Y(n1986) );
  MUX2X1 U6027 ( .B(n1990), .A(n1991), .S(n3083), .Y(n1989) );
  MUX2X1 U6028 ( .B(n1993), .A(n1994), .S(n3083), .Y(n1992) );
  MUX2X1 U6029 ( .B(n1996), .A(n1997), .S(n3083), .Y(n1995) );
  MUX2X1 U6030 ( .B(n1999), .A(n2000), .S(n3083), .Y(n1998) );
  MUX2X1 U6031 ( .B(n2002), .A(n2003), .S(n3175), .Y(n2001) );
  MUX2X1 U6032 ( .B(n2004), .A(n2005), .S(n18), .Y(data_out[26]) );
  MUX2X1 U6033 ( .B(n2007), .A(n2008), .S(n3083), .Y(n2006) );
  MUX2X1 U6034 ( .B(n2010), .A(n2011), .S(n3083), .Y(n2009) );
  MUX2X1 U6035 ( .B(n2013), .A(n2014), .S(n3083), .Y(n2012) );
  MUX2X1 U6036 ( .B(n2016), .A(n2017), .S(n3083), .Y(n2015) );
  MUX2X1 U6037 ( .B(n2019), .A(n2020), .S(n3175), .Y(n2018) );
  MUX2X1 U6038 ( .B(n2022), .A(n2023), .S(n3083), .Y(n2021) );
  MUX2X1 U6039 ( .B(n2025), .A(n2026), .S(n3083), .Y(n2024) );
  MUX2X1 U6040 ( .B(n2028), .A(n2029), .S(n3083), .Y(n2027) );
  MUX2X1 U6041 ( .B(n2031), .A(n2032), .S(n3083), .Y(n2030) );
  MUX2X1 U6042 ( .B(n2034), .A(n2035), .S(n3175), .Y(n2033) );
  MUX2X1 U6043 ( .B(n2037), .A(n2038), .S(n3084), .Y(n2036) );
  MUX2X1 U6044 ( .B(n2040), .A(n2041), .S(n3084), .Y(n2039) );
  MUX2X1 U6045 ( .B(n2043), .A(n2044), .S(n3084), .Y(n2042) );
  MUX2X1 U6046 ( .B(n2046), .A(n2047), .S(n3084), .Y(n2045) );
  MUX2X1 U6047 ( .B(n2049), .A(n2050), .S(n3175), .Y(n2048) );
  MUX2X1 U6048 ( .B(n2052), .A(n2053), .S(n3084), .Y(n2051) );
  MUX2X1 U6049 ( .B(n2055), .A(n2056), .S(n3084), .Y(n2054) );
  MUX2X1 U6050 ( .B(n2058), .A(n2059), .S(n3084), .Y(n2057) );
  MUX2X1 U6051 ( .B(n2061), .A(n2062), .S(n3084), .Y(n2060) );
  MUX2X1 U6052 ( .B(n2064), .A(n2065), .S(n3175), .Y(n2063) );
  MUX2X1 U6053 ( .B(n2066), .A(n2067), .S(n18), .Y(data_out[27]) );
  MUX2X1 U6054 ( .B(n2069), .A(n2070), .S(n3084), .Y(n2068) );
  MUX2X1 U6055 ( .B(n2072), .A(n2073), .S(n3084), .Y(n2071) );
  MUX2X1 U6056 ( .B(n2075), .A(n2076), .S(n3084), .Y(n2074) );
  MUX2X1 U6057 ( .B(n2078), .A(n2079), .S(n3084), .Y(n2077) );
  MUX2X1 U6058 ( .B(n2081), .A(n2082), .S(n3175), .Y(n2080) );
  MUX2X1 U6059 ( .B(n2084), .A(n2085), .S(n3085), .Y(n2083) );
  MUX2X1 U6060 ( .B(n2087), .A(n2088), .S(n3085), .Y(n2086) );
  MUX2X1 U6061 ( .B(n2090), .A(n2091), .S(n3085), .Y(n2089) );
  MUX2X1 U6062 ( .B(n2093), .A(n2094), .S(n3085), .Y(n2092) );
  MUX2X1 U6063 ( .B(n2096), .A(n2097), .S(n3175), .Y(n2095) );
  MUX2X1 U6064 ( .B(n2099), .A(n2100), .S(n3085), .Y(n2098) );
  MUX2X1 U6065 ( .B(n2102), .A(n2103), .S(n3085), .Y(n2101) );
  MUX2X1 U6066 ( .B(n2105), .A(n2106), .S(n3085), .Y(n2104) );
  MUX2X1 U6067 ( .B(n2108), .A(n2109), .S(n3085), .Y(n2107) );
  MUX2X1 U6068 ( .B(n2111), .A(n2112), .S(n3175), .Y(n2110) );
  MUX2X1 U6069 ( .B(n2114), .A(n2115), .S(n3085), .Y(n2113) );
  MUX2X1 U6070 ( .B(n2117), .A(n2118), .S(n3085), .Y(n2116) );
  MUX2X1 U6071 ( .B(n2120), .A(n2121), .S(n3085), .Y(n2119) );
  MUX2X1 U6072 ( .B(n2123), .A(n2124), .S(n3085), .Y(n2122) );
  MUX2X1 U6073 ( .B(n2126), .A(n2127), .S(n3175), .Y(n2125) );
  MUX2X1 U6074 ( .B(n2128), .A(n2129), .S(n18), .Y(data_out[28]) );
  MUX2X1 U6075 ( .B(n2131), .A(n2132), .S(n3086), .Y(n2130) );
  MUX2X1 U6076 ( .B(n2134), .A(n2135), .S(n3086), .Y(n2133) );
  MUX2X1 U6077 ( .B(n2137), .A(n2138), .S(n3086), .Y(n2136) );
  MUX2X1 U6078 ( .B(n2140), .A(n2141), .S(n3086), .Y(n2139) );
  MUX2X1 U6079 ( .B(n2143), .A(n2144), .S(n3176), .Y(n2142) );
  MUX2X1 U6080 ( .B(n2146), .A(n2147), .S(n3086), .Y(n2145) );
  MUX2X1 U6081 ( .B(n2149), .A(n2150), .S(n3086), .Y(n2148) );
  MUX2X1 U6082 ( .B(n2152), .A(n2153), .S(n3086), .Y(n2151) );
  MUX2X1 U6083 ( .B(n2155), .A(n2156), .S(n3086), .Y(n2154) );
  MUX2X1 U6084 ( .B(n2158), .A(n2159), .S(n3176), .Y(n2157) );
  MUX2X1 U6085 ( .B(n2161), .A(n2162), .S(n3086), .Y(n2160) );
  MUX2X1 U6086 ( .B(n2164), .A(n2165), .S(n3086), .Y(n2163) );
  MUX2X1 U6087 ( .B(n2167), .A(n2168), .S(n3086), .Y(n2166) );
  MUX2X1 U6088 ( .B(n2170), .A(n2171), .S(n3086), .Y(n2169) );
  MUX2X1 U6089 ( .B(n2173), .A(n2174), .S(n3176), .Y(n2172) );
  MUX2X1 U6090 ( .B(n2176), .A(n2177), .S(n3087), .Y(n2175) );
  MUX2X1 U6091 ( .B(n2179), .A(n2180), .S(n3087), .Y(n2178) );
  MUX2X1 U6092 ( .B(n2182), .A(n2183), .S(n3087), .Y(n2181) );
  MUX2X1 U6093 ( .B(n2185), .A(n2186), .S(n3087), .Y(n2184) );
  MUX2X1 U6094 ( .B(n2188), .A(n2189), .S(n3176), .Y(n2187) );
  MUX2X1 U6095 ( .B(n2190), .A(n2191), .S(n18), .Y(data_out[29]) );
  MUX2X1 U6096 ( .B(n2193), .A(n2194), .S(n3087), .Y(n2192) );
  MUX2X1 U6097 ( .B(n2196), .A(n2197), .S(n3087), .Y(n2195) );
  MUX2X1 U6098 ( .B(n2199), .A(n2200), .S(n3087), .Y(n2198) );
  MUX2X1 U6099 ( .B(n2202), .A(n2203), .S(n3087), .Y(n2201) );
  MUX2X1 U6100 ( .B(n2205), .A(n2206), .S(n3176), .Y(n2204) );
  MUX2X1 U6101 ( .B(n2208), .A(n2209), .S(n3087), .Y(n2207) );
  MUX2X1 U6102 ( .B(n2211), .A(n2212), .S(n3087), .Y(n2210) );
  MUX2X1 U6103 ( .B(n2214), .A(n2215), .S(n3087), .Y(n2213) );
  MUX2X1 U6104 ( .B(n2217), .A(n2218), .S(n3087), .Y(n2216) );
  MUX2X1 U6105 ( .B(n2220), .A(n2221), .S(n3176), .Y(n2219) );
  MUX2X1 U6106 ( .B(n2223), .A(n2224), .S(n3088), .Y(n2222) );
  MUX2X1 U6107 ( .B(n2226), .A(n2227), .S(n3088), .Y(n2225) );
  MUX2X1 U6108 ( .B(n2229), .A(n2230), .S(n3088), .Y(n2228) );
  MUX2X1 U6109 ( .B(n2232), .A(n2233), .S(n3088), .Y(n2231) );
  MUX2X1 U6110 ( .B(n2235), .A(n2236), .S(n3176), .Y(n2234) );
  MUX2X1 U6111 ( .B(n2238), .A(n2239), .S(n3088), .Y(n2237) );
  MUX2X1 U6112 ( .B(n2241), .A(n2242), .S(n3088), .Y(n2240) );
  MUX2X1 U6113 ( .B(n2244), .A(n2245), .S(n3088), .Y(n2243) );
  MUX2X1 U6114 ( .B(n2247), .A(n2248), .S(n3088), .Y(n2246) );
  MUX2X1 U6115 ( .B(n2250), .A(n2251), .S(n3176), .Y(n2249) );
  MUX2X1 U6116 ( .B(n2252), .A(n2253), .S(n18), .Y(data_out[30]) );
  MUX2X1 U6117 ( .B(n2255), .A(n2256), .S(n3088), .Y(n2254) );
  MUX2X1 U6118 ( .B(n2258), .A(n2259), .S(n3088), .Y(n2257) );
  MUX2X1 U6119 ( .B(n2261), .A(n2262), .S(n3088), .Y(n2260) );
  MUX2X1 U6120 ( .B(n2264), .A(n2265), .S(n3088), .Y(n2263) );
  MUX2X1 U6121 ( .B(n2267), .A(n2268), .S(n3176), .Y(n2266) );
  MUX2X1 U6122 ( .B(n2270), .A(n2271), .S(n3089), .Y(n2269) );
  MUX2X1 U6123 ( .B(n2273), .A(n2274), .S(n3089), .Y(n2272) );
  MUX2X1 U6124 ( .B(n2276), .A(n2277), .S(n3089), .Y(n2275) );
  MUX2X1 U6125 ( .B(n2279), .A(n2280), .S(n3089), .Y(n2278) );
  MUX2X1 U6126 ( .B(n2282), .A(n2283), .S(n3176), .Y(n2281) );
  MUX2X1 U6127 ( .B(n2285), .A(n2286), .S(n3089), .Y(n2284) );
  MUX2X1 U6128 ( .B(n2288), .A(n2289), .S(n3089), .Y(n2287) );
  MUX2X1 U6129 ( .B(n2291), .A(n2292), .S(n3089), .Y(n2290) );
  MUX2X1 U6130 ( .B(n2294), .A(n2295), .S(n3089), .Y(n2293) );
  MUX2X1 U6131 ( .B(n2297), .A(n2298), .S(n3176), .Y(n2296) );
  MUX2X1 U6132 ( .B(n2300), .A(n2301), .S(n3089), .Y(n2299) );
  MUX2X1 U6133 ( .B(n2303), .A(n2304), .S(n3089), .Y(n2302) );
  MUX2X1 U6134 ( .B(n2306), .A(n2307), .S(n3089), .Y(n2305) );
  MUX2X1 U6135 ( .B(n2309), .A(n2310), .S(n3089), .Y(n2308) );
  MUX2X1 U6136 ( .B(n2312), .A(n2313), .S(n3176), .Y(n2311) );
  MUX2X1 U6137 ( .B(n2314), .A(n2315), .S(n18), .Y(data_out[31]) );
  MUX2X1 U6138 ( .B(n2317), .A(n2318), .S(n3090), .Y(n2316) );
  MUX2X1 U6139 ( .B(n2320), .A(n2321), .S(n3090), .Y(n2319) );
  MUX2X1 U6140 ( .B(n2323), .A(n2324), .S(n3090), .Y(n2322) );
  MUX2X1 U6141 ( .B(n2326), .A(n2327), .S(n3090), .Y(n2325) );
  MUX2X1 U6142 ( .B(n2329), .A(n2330), .S(n3177), .Y(n2328) );
  MUX2X1 U6143 ( .B(n2332), .A(n2333), .S(n3090), .Y(n2331) );
  MUX2X1 U6144 ( .B(n2335), .A(n2336), .S(n3090), .Y(n2334) );
  MUX2X1 U6145 ( .B(n2338), .A(n2339), .S(n3090), .Y(n2337) );
  MUX2X1 U6146 ( .B(n2341), .A(n2342), .S(n3090), .Y(n2340) );
  MUX2X1 U6147 ( .B(n2344), .A(n2345), .S(n3177), .Y(n2343) );
  MUX2X1 U6148 ( .B(n2347), .A(n2348), .S(n3090), .Y(n2346) );
  MUX2X1 U6149 ( .B(n2350), .A(n2351), .S(n3090), .Y(n2349) );
  MUX2X1 U6150 ( .B(n2353), .A(n2354), .S(n3090), .Y(n2352) );
  MUX2X1 U6151 ( .B(n2356), .A(n2357), .S(n3090), .Y(n2355) );
  MUX2X1 U6152 ( .B(n2359), .A(n2360), .S(n3177), .Y(n2358) );
  MUX2X1 U6153 ( .B(n2362), .A(n2363), .S(n3091), .Y(n2361) );
  MUX2X1 U6154 ( .B(n2365), .A(n2366), .S(n3091), .Y(n2364) );
  MUX2X1 U6155 ( .B(n2368), .A(n2369), .S(n3091), .Y(n2367) );
  MUX2X1 U6156 ( .B(n2371), .A(n2372), .S(n3091), .Y(n2370) );
  MUX2X1 U6157 ( .B(n2374), .A(n2375), .S(n3177), .Y(n2373) );
  MUX2X1 U6158 ( .B(n2376), .A(n2377), .S(n18), .Y(data_out[32]) );
  MUX2X1 U6159 ( .B(n2379), .A(n2380), .S(n3091), .Y(n2378) );
  MUX2X1 U6160 ( .B(n2382), .A(n2383), .S(n3091), .Y(n2381) );
  MUX2X1 U6161 ( .B(n2385), .A(n2386), .S(n3091), .Y(n2384) );
  MUX2X1 U6162 ( .B(n2388), .A(n2389), .S(n3091), .Y(n2387) );
  MUX2X1 U6163 ( .B(n2391), .A(n2392), .S(n3177), .Y(n2390) );
  MUX2X1 U6164 ( .B(n2394), .A(n2395), .S(n3091), .Y(n2393) );
  MUX2X1 U6165 ( .B(n2397), .A(n2398), .S(n3091), .Y(n2396) );
  MUX2X1 U6166 ( .B(n2400), .A(n2401), .S(n3091), .Y(n2399) );
  MUX2X1 U6167 ( .B(n2403), .A(n2404), .S(n3091), .Y(n2402) );
  MUX2X1 U6168 ( .B(n2406), .A(n2407), .S(n3177), .Y(n2405) );
  MUX2X1 U6169 ( .B(n2409), .A(n2410), .S(n3092), .Y(n2408) );
  MUX2X1 U6170 ( .B(n2412), .A(n2413), .S(n3092), .Y(n2411) );
  MUX2X1 U6171 ( .B(n2415), .A(n2416), .S(n3092), .Y(n2414) );
  MUX2X1 U6172 ( .B(n2418), .A(n2419), .S(n3092), .Y(n2417) );
  MUX2X1 U6173 ( .B(n2421), .A(n2422), .S(n3177), .Y(n2420) );
  MUX2X1 U6174 ( .B(n2424), .A(n2425), .S(n3092), .Y(n2423) );
  MUX2X1 U6175 ( .B(n2427), .A(n2428), .S(n3092), .Y(n2426) );
  MUX2X1 U6176 ( .B(n2430), .A(n2431), .S(n3092), .Y(n2429) );
  MUX2X1 U6177 ( .B(n2433), .A(n2434), .S(n3092), .Y(n2432) );
  MUX2X1 U6178 ( .B(n2436), .A(n2437), .S(n3177), .Y(n2435) );
  MUX2X1 U6179 ( .B(n2438), .A(n2439), .S(n18), .Y(data_out[33]) );
  MUX2X1 U6180 ( .B(n2441), .A(n2442), .S(n3092), .Y(n2440) );
  MUX2X1 U6181 ( .B(n2444), .A(n2445), .S(n3092), .Y(n2443) );
  MUX2X1 U6182 ( .B(n2447), .A(n2448), .S(n3092), .Y(n2446) );
  MUX2X1 U6183 ( .B(n2450), .A(n2451), .S(n3092), .Y(n2449) );
  MUX2X1 U6184 ( .B(n2453), .A(n2454), .S(n3177), .Y(n2452) );
  MUX2X1 U6185 ( .B(n2456), .A(n2457), .S(n3093), .Y(n2455) );
  MUX2X1 U6186 ( .B(n2459), .A(n2460), .S(n3093), .Y(n2458) );
  MUX2X1 U6187 ( .B(n2462), .A(n2463), .S(n3093), .Y(n2461) );
  MUX2X1 U6188 ( .B(n2465), .A(n2466), .S(n3093), .Y(n2464) );
  MUX2X1 U6189 ( .B(n2468), .A(n2469), .S(n3177), .Y(n2467) );
  MUX2X1 U6190 ( .B(n2471), .A(n2472), .S(n3093), .Y(n2470) );
  MUX2X1 U6191 ( .B(n2474), .A(n2475), .S(n3093), .Y(n2473) );
  MUX2X1 U6192 ( .B(n2477), .A(n2478), .S(n3093), .Y(n2476) );
  MUX2X1 U6193 ( .B(n2480), .A(n2481), .S(n3093), .Y(n2479) );
  MUX2X1 U6194 ( .B(n2483), .A(n2484), .S(n3177), .Y(n2482) );
  MUX2X1 U6195 ( .B(n2486), .A(n2487), .S(n3093), .Y(n2485) );
  MUX2X1 U6196 ( .B(n2489), .A(n2490), .S(n3093), .Y(n2488) );
  MUX2X1 U6197 ( .B(n2492), .A(n2493), .S(n3093), .Y(n2491) );
  MUX2X1 U6198 ( .B(n2495), .A(n2496), .S(n3093), .Y(n2494) );
  MUX2X1 U6199 ( .B(n2498), .A(n2499), .S(n3177), .Y(n2497) );
  MUX2X1 U6200 ( .B(n2500), .A(n2501), .S(n18), .Y(data_out[34]) );
  MUX2X1 U6201 ( .B(n2503), .A(n2504), .S(n3094), .Y(n2502) );
  MUX2X1 U6202 ( .B(n2506), .A(n2507), .S(n3094), .Y(n2505) );
  MUX2X1 U6203 ( .B(n2509), .A(n2510), .S(n3094), .Y(n2508) );
  MUX2X1 U6204 ( .B(n2512), .A(n2513), .S(n3094), .Y(n2511) );
  MUX2X1 U6205 ( .B(n2515), .A(n2516), .S(n3178), .Y(n2514) );
  MUX2X1 U6206 ( .B(n2518), .A(n2519), .S(n3094), .Y(n2517) );
  MUX2X1 U6207 ( .B(n2521), .A(n2522), .S(n3094), .Y(n2520) );
  MUX2X1 U6208 ( .B(n2524), .A(n2525), .S(n3094), .Y(n2523) );
  MUX2X1 U6209 ( .B(n2527), .A(n2528), .S(n3094), .Y(n2526) );
  MUX2X1 U6210 ( .B(n2530), .A(n2531), .S(n3178), .Y(n2529) );
  MUX2X1 U6211 ( .B(n2533), .A(n2534), .S(n3094), .Y(n2532) );
  MUX2X1 U6212 ( .B(n2536), .A(n2537), .S(n3094), .Y(n2535) );
  MUX2X1 U6213 ( .B(n2539), .A(n2540), .S(n3094), .Y(n2538) );
  MUX2X1 U6214 ( .B(n2542), .A(n2543), .S(n3094), .Y(n2541) );
  MUX2X1 U6215 ( .B(n2545), .A(n2546), .S(n3178), .Y(n2544) );
  MUX2X1 U6216 ( .B(n2548), .A(n2549), .S(n3095), .Y(n2547) );
  MUX2X1 U6217 ( .B(n2551), .A(n2552), .S(n3095), .Y(n2550) );
  MUX2X1 U6218 ( .B(n2554), .A(n2555), .S(n3095), .Y(n2553) );
  MUX2X1 U6219 ( .B(n2557), .A(n2558), .S(n3095), .Y(n2556) );
  MUX2X1 U6220 ( .B(n2560), .A(n2561), .S(n3178), .Y(n2559) );
  MUX2X1 U6221 ( .B(n2562), .A(n2563), .S(n18), .Y(data_out[35]) );
  MUX2X1 U6222 ( .B(n2565), .A(n2566), .S(n3095), .Y(n2564) );
  MUX2X1 U6223 ( .B(n2568), .A(n2569), .S(n3095), .Y(n2567) );
  MUX2X1 U6224 ( .B(n2571), .A(n2572), .S(n3095), .Y(n2570) );
  MUX2X1 U6225 ( .B(n2574), .A(n2575), .S(n3095), .Y(n2573) );
  MUX2X1 U6226 ( .B(n2577), .A(n2578), .S(n3178), .Y(n2576) );
  MUX2X1 U6227 ( .B(n2580), .A(n2581), .S(n3095), .Y(n2579) );
  MUX2X1 U6228 ( .B(n2583), .A(n2584), .S(n3095), .Y(n2582) );
  MUX2X1 U6229 ( .B(n2586), .A(n2587), .S(n3095), .Y(n2585) );
  MUX2X1 U6230 ( .B(n2589), .A(n2590), .S(n3095), .Y(n2588) );
  MUX2X1 U6231 ( .B(n2592), .A(n2593), .S(n3178), .Y(n2591) );
  MUX2X1 U6232 ( .B(n2595), .A(n2596), .S(n3096), .Y(n2594) );
  MUX2X1 U6233 ( .B(n2598), .A(n2599), .S(n3096), .Y(n2597) );
  MUX2X1 U6234 ( .B(n2601), .A(n2602), .S(n3096), .Y(n2600) );
  MUX2X1 U6235 ( .B(n2604), .A(n2605), .S(n3096), .Y(n2603) );
  MUX2X1 U6236 ( .B(n2607), .A(n2608), .S(n3178), .Y(n2606) );
  MUX2X1 U6237 ( .B(n2610), .A(n2611), .S(n3096), .Y(n2609) );
  MUX2X1 U6238 ( .B(n2613), .A(n2614), .S(n3096), .Y(n2612) );
  MUX2X1 U6239 ( .B(n2616), .A(n2617), .S(n3096), .Y(n2615) );
  MUX2X1 U6240 ( .B(n2619), .A(n2620), .S(n3096), .Y(n2618) );
  MUX2X1 U6241 ( .B(n2622), .A(n2623), .S(n3178), .Y(n2621) );
  MUX2X1 U6242 ( .B(n2624), .A(n2625), .S(n18), .Y(data_out[36]) );
  MUX2X1 U6243 ( .B(n2627), .A(n2628), .S(n3096), .Y(n2626) );
  MUX2X1 U6244 ( .B(n2630), .A(n2631), .S(n3096), .Y(n2629) );
  MUX2X1 U6245 ( .B(n2633), .A(n2634), .S(n3096), .Y(n2632) );
  MUX2X1 U6246 ( .B(n2636), .A(n2637), .S(n3096), .Y(n2635) );
  MUX2X1 U6247 ( .B(n2639), .A(n2640), .S(n3178), .Y(n2638) );
  MUX2X1 U6248 ( .B(n2642), .A(n2643), .S(n3097), .Y(n2641) );
  MUX2X1 U6249 ( .B(n2645), .A(n2646), .S(n3097), .Y(n2644) );
  MUX2X1 U6250 ( .B(n2648), .A(n2649), .S(n3097), .Y(n2647) );
  MUX2X1 U6251 ( .B(n2651), .A(n2652), .S(n3097), .Y(n2650) );
  MUX2X1 U6252 ( .B(n2654), .A(n2655), .S(n3178), .Y(n2653) );
  MUX2X1 U6253 ( .B(n2657), .A(n2658), .S(n3097), .Y(n2656) );
  MUX2X1 U6254 ( .B(n2660), .A(n2661), .S(n3097), .Y(n2659) );
  MUX2X1 U6255 ( .B(n2663), .A(n2664), .S(n3097), .Y(n2662) );
  MUX2X1 U6256 ( .B(n2666), .A(n2667), .S(n3097), .Y(n2665) );
  MUX2X1 U6257 ( .B(n2669), .A(n2670), .S(n3178), .Y(n2668) );
  MUX2X1 U6258 ( .B(n2672), .A(n2673), .S(n3097), .Y(n2671) );
  MUX2X1 U6259 ( .B(n2675), .A(n2676), .S(n3097), .Y(n2674) );
  MUX2X1 U6260 ( .B(n2678), .A(n2679), .S(n3097), .Y(n2677) );
  MUX2X1 U6261 ( .B(n2681), .A(n2682), .S(n3097), .Y(n2680) );
  MUX2X1 U6262 ( .B(n2684), .A(n2685), .S(n3178), .Y(n2683) );
  MUX2X1 U6263 ( .B(n2686), .A(n2687), .S(n18), .Y(data_out[37]) );
  MUX2X1 U6264 ( .B(n2689), .A(n2690), .S(n3098), .Y(n2688) );
  MUX2X1 U6265 ( .B(n2692), .A(n2693), .S(n3098), .Y(n2691) );
  MUX2X1 U6266 ( .B(n2695), .A(n2696), .S(n3098), .Y(n2694) );
  MUX2X1 U6267 ( .B(n2698), .A(n2699), .S(n3098), .Y(n2697) );
  MUX2X1 U6268 ( .B(n2701), .A(n2702), .S(n3179), .Y(n2700) );
  MUX2X1 U6269 ( .B(n2704), .A(n2705), .S(n3098), .Y(n2703) );
  MUX2X1 U6270 ( .B(n2707), .A(n2708), .S(n3098), .Y(n2706) );
  MUX2X1 U6271 ( .B(n2710), .A(n2711), .S(n3098), .Y(n2709) );
  MUX2X1 U6272 ( .B(n2713), .A(n2714), .S(n3098), .Y(n2712) );
  MUX2X1 U6273 ( .B(n2716), .A(n2717), .S(n3179), .Y(n2715) );
  MUX2X1 U6274 ( .B(n2719), .A(n2720), .S(n3098), .Y(n2718) );
  MUX2X1 U6275 ( .B(n2722), .A(n2723), .S(n3098), .Y(n2721) );
  MUX2X1 U6276 ( .B(n2738), .A(n2739), .S(n3098), .Y(n2724) );
  MUX2X1 U6277 ( .B(n2741), .A(n2742), .S(n3098), .Y(n2740) );
  MUX2X1 U6278 ( .B(n2744), .A(n2745), .S(n3179), .Y(n2743) );
  MUX2X1 U6279 ( .B(n2747), .A(n2748), .S(n3099), .Y(n2746) );
  MUX2X1 U6280 ( .B(n2750), .A(n2751), .S(n3099), .Y(n2749) );
  MUX2X1 U6281 ( .B(n2753), .A(n2754), .S(n3099), .Y(n2752) );
  MUX2X1 U6282 ( .B(n2756), .A(n2757), .S(n3099), .Y(n2755) );
  MUX2X1 U6283 ( .B(n2759), .A(n2760), .S(n3179), .Y(n2758) );
  MUX2X1 U6284 ( .B(n2761), .A(n2762), .S(n18), .Y(data_out[38]) );
  MUX2X1 U6285 ( .B(n2764), .A(n2765), .S(n3099), .Y(n2763) );
  MUX2X1 U6286 ( .B(n2767), .A(n2768), .S(n3099), .Y(n2766) );
  MUX2X1 U6287 ( .B(n2770), .A(n2771), .S(n3099), .Y(n2769) );
  MUX2X1 U6288 ( .B(n2773), .A(n2774), .S(n3099), .Y(n2772) );
  MUX2X1 U6289 ( .B(n2776), .A(n2777), .S(n3179), .Y(n2775) );
  MUX2X1 U6290 ( .B(n2779), .A(n2780), .S(n3099), .Y(n2778) );
  MUX2X1 U6291 ( .B(n2782), .A(n2783), .S(n3099), .Y(n2781) );
  MUX2X1 U6292 ( .B(n2785), .A(n2786), .S(n3099), .Y(n2784) );
  MUX2X1 U6293 ( .B(n2788), .A(n2789), .S(n3099), .Y(n2787) );
  MUX2X1 U6294 ( .B(n2791), .A(n2792), .S(n3179), .Y(n2790) );
  MUX2X1 U6295 ( .B(n2794), .A(n2795), .S(n3100), .Y(n2793) );
  MUX2X1 U6296 ( .B(n2797), .A(n2798), .S(n3100), .Y(n2796) );
  MUX2X1 U6297 ( .B(n2800), .A(n2801), .S(n3100), .Y(n2799) );
  MUX2X1 U6298 ( .B(n2803), .A(n2804), .S(n3100), .Y(n2802) );
  MUX2X1 U6299 ( .B(n2806), .A(n2807), .S(n3179), .Y(n2805) );
  MUX2X1 U6300 ( .B(n2809), .A(n2810), .S(n3100), .Y(n2808) );
  MUX2X1 U6301 ( .B(n2812), .A(n2813), .S(n3100), .Y(n2811) );
  MUX2X1 U6302 ( .B(n2815), .A(n2816), .S(n3100), .Y(n2814) );
  MUX2X1 U6303 ( .B(n2818), .A(n2819), .S(n3100), .Y(n2817) );
  MUX2X1 U6304 ( .B(n2821), .A(n2822), .S(n3179), .Y(n2820) );
  MUX2X1 U6305 ( .B(n2823), .A(n2824), .S(n18), .Y(data_out[39]) );
  MUX2X1 U6306 ( .B(n2826), .A(n2827), .S(n3100), .Y(n2825) );
  MUX2X1 U6307 ( .B(n2829), .A(n2830), .S(n3100), .Y(n2828) );
  MUX2X1 U6308 ( .B(n2832), .A(n2833), .S(n3100), .Y(n2831) );
  MUX2X1 U6309 ( .B(n2835), .A(n2836), .S(n3100), .Y(n2834) );
  MUX2X1 U6310 ( .B(n2838), .A(n2839), .S(n3179), .Y(n2837) );
  MUX2X1 U6311 ( .B(n2841), .A(n2842), .S(n3101), .Y(n2840) );
  MUX2X1 U6312 ( .B(n2844), .A(n2845), .S(n3101), .Y(n2843) );
  MUX2X1 U6313 ( .B(n2847), .A(n2848), .S(n3101), .Y(n2846) );
  MUX2X1 U6314 ( .B(n2850), .A(n2851), .S(n3101), .Y(n2849) );
  MUX2X1 U6315 ( .B(n2853), .A(n2854), .S(n3179), .Y(n2852) );
  MUX2X1 U6316 ( .B(n2856), .A(n2857), .S(n3101), .Y(n2855) );
  MUX2X1 U6317 ( .B(n2859), .A(n2860), .S(n3101), .Y(n2858) );
  MUX2X1 U6318 ( .B(n2862), .A(n2863), .S(n3101), .Y(n2861) );
  MUX2X1 U6319 ( .B(n2865), .A(n2866), .S(n3101), .Y(n2864) );
  MUX2X1 U6320 ( .B(n2868), .A(n2869), .S(n3179), .Y(n2867) );
  MUX2X1 U6321 ( .B(n2871), .A(n2872), .S(n3101), .Y(n2870) );
  MUX2X1 U6322 ( .B(n2874), .A(n2875), .S(n3101), .Y(n2873) );
  MUX2X1 U6323 ( .B(n2877), .A(n2878), .S(n3101), .Y(n2876) );
  MUX2X1 U6324 ( .B(n2880), .A(n2881), .S(n3101), .Y(n2879) );
  MUX2X1 U6325 ( .B(n2883), .A(n2884), .S(n3179), .Y(n2882) );
  MUX2X1 U6326 ( .B(n2885), .A(n2886), .S(n18), .Y(data_out[40]) );
  MUX2X1 U6327 ( .B(arr[2542]), .A(arr[2583]), .S(n2924), .Y(n334) );
  MUX2X1 U6328 ( .B(arr[2460]), .A(arr[2501]), .S(n2924), .Y(n333) );
  MUX2X1 U6329 ( .B(arr[2378]), .A(arr[2419]), .S(n2924), .Y(n337) );
  MUX2X1 U6330 ( .B(arr[2296]), .A(arr[2337]), .S(n2924), .Y(n336) );
  MUX2X1 U6331 ( .B(n335), .A(n332), .S(n3128), .Y(n346) );
  MUX2X1 U6332 ( .B(arr[2214]), .A(arr[2255]), .S(n2925), .Y(n340) );
  MUX2X1 U6333 ( .B(arr[2132]), .A(arr[2173]), .S(n2925), .Y(n339) );
  MUX2X1 U6334 ( .B(arr[2050]), .A(arr[2091]), .S(n2925), .Y(n343) );
  MUX2X1 U6335 ( .B(arr[1968]), .A(arr[2009]), .S(n2925), .Y(n342) );
  MUX2X1 U6336 ( .B(n341), .A(n338), .S(n3128), .Y(n345) );
  MUX2X1 U6337 ( .B(arr[1886]), .A(arr[1927]), .S(n2925), .Y(n349) );
  MUX2X1 U6338 ( .B(arr[1804]), .A(arr[1845]), .S(n2925), .Y(n348) );
  MUX2X1 U6339 ( .B(arr[1722]), .A(arr[1763]), .S(n2925), .Y(n352) );
  MUX2X1 U6340 ( .B(arr[1640]), .A(arr[1681]), .S(n2925), .Y(n351) );
  MUX2X1 U6341 ( .B(n350), .A(n347), .S(n3128), .Y(n361) );
  MUX2X1 U6342 ( .B(arr[1558]), .A(arr[1599]), .S(n2925), .Y(n355) );
  MUX2X1 U6343 ( .B(arr[1476]), .A(arr[1517]), .S(n2925), .Y(n354) );
  MUX2X1 U6344 ( .B(arr[1394]), .A(arr[1435]), .S(n2925), .Y(n358) );
  MUX2X1 U6345 ( .B(arr[1312]), .A(arr[1353]), .S(n2925), .Y(n357) );
  MUX2X1 U6346 ( .B(n356), .A(n353), .S(n3128), .Y(n360) );
  MUX2X1 U6347 ( .B(n359), .A(n344), .S(n3180), .Y(n393) );
  MUX2X1 U6348 ( .B(arr[1230]), .A(arr[1271]), .S(n2926), .Y(n364) );
  MUX2X1 U6349 ( .B(arr[1148]), .A(arr[1189]), .S(n2926), .Y(n363) );
  MUX2X1 U6350 ( .B(arr[1066]), .A(arr[1107]), .S(n2926), .Y(n367) );
  MUX2X1 U6351 ( .B(arr[984]), .A(arr[1025]), .S(n2926), .Y(n366) );
  MUX2X1 U6352 ( .B(n365), .A(n362), .S(n3129), .Y(n376) );
  MUX2X1 U6353 ( .B(arr[902]), .A(arr[943]), .S(n2926), .Y(n370) );
  MUX2X1 U6354 ( .B(arr[820]), .A(arr[861]), .S(n2926), .Y(n369) );
  MUX2X1 U6355 ( .B(arr[738]), .A(arr[779]), .S(n2926), .Y(n373) );
  MUX2X1 U6356 ( .B(arr[656]), .A(arr[697]), .S(n2926), .Y(n372) );
  MUX2X1 U6357 ( .B(n371), .A(n368), .S(n3129), .Y(n375) );
  MUX2X1 U6358 ( .B(arr[574]), .A(arr[615]), .S(n2926), .Y(n379) );
  MUX2X1 U6359 ( .B(arr[492]), .A(arr[533]), .S(n2926), .Y(n378) );
  MUX2X1 U6360 ( .B(arr[410]), .A(arr[451]), .S(n2926), .Y(n382) );
  MUX2X1 U6361 ( .B(arr[328]), .A(arr[369]), .S(n2926), .Y(n381) );
  MUX2X1 U6362 ( .B(n380), .A(n377), .S(n3129), .Y(n391) );
  MUX2X1 U6363 ( .B(arr[246]), .A(arr[287]), .S(n2927), .Y(n385) );
  MUX2X1 U6364 ( .B(arr[164]), .A(arr[205]), .S(n2927), .Y(n384) );
  MUX2X1 U6365 ( .B(arr[82]), .A(arr[123]), .S(n2927), .Y(n388) );
  MUX2X1 U6366 ( .B(arr[0]), .A(arr[41]), .S(n2927), .Y(n387) );
  MUX2X1 U6367 ( .B(n386), .A(n383), .S(n3129), .Y(n390) );
  MUX2X1 U6368 ( .B(n389), .A(n374), .S(n3180), .Y(n392) );
  MUX2X1 U6369 ( .B(arr[2543]), .A(arr[2584]), .S(n2927), .Y(n396) );
  MUX2X1 U6370 ( .B(arr[2461]), .A(arr[2502]), .S(n2927), .Y(n395) );
  MUX2X1 U6371 ( .B(arr[2379]), .A(arr[2420]), .S(n2927), .Y(n399) );
  MUX2X1 U6372 ( .B(arr[2297]), .A(arr[2338]), .S(n2927), .Y(n398) );
  MUX2X1 U6373 ( .B(n397), .A(n394), .S(n3129), .Y(n408) );
  MUX2X1 U6374 ( .B(arr[2215]), .A(arr[2256]), .S(n2927), .Y(n402) );
  MUX2X1 U6375 ( .B(arr[2133]), .A(arr[2174]), .S(n2927), .Y(n401) );
  MUX2X1 U6376 ( .B(arr[2051]), .A(arr[2092]), .S(n2927), .Y(n405) );
  MUX2X1 U6377 ( .B(arr[1969]), .A(arr[2010]), .S(n2927), .Y(n404) );
  MUX2X1 U6378 ( .B(n403), .A(n400), .S(n3129), .Y(n407) );
  MUX2X1 U6379 ( .B(arr[1887]), .A(arr[1928]), .S(n2928), .Y(n411) );
  MUX2X1 U6380 ( .B(arr[1805]), .A(arr[1846]), .S(n2928), .Y(n410) );
  MUX2X1 U6381 ( .B(arr[1723]), .A(arr[1764]), .S(n2928), .Y(n414) );
  MUX2X1 U6382 ( .B(arr[1641]), .A(arr[1682]), .S(n2928), .Y(n413) );
  MUX2X1 U6383 ( .B(n412), .A(n409), .S(n3129), .Y(n423) );
  MUX2X1 U6384 ( .B(arr[1559]), .A(arr[1600]), .S(n2928), .Y(n417) );
  MUX2X1 U6385 ( .B(arr[1477]), .A(arr[1518]), .S(n2928), .Y(n416) );
  MUX2X1 U6386 ( .B(arr[1395]), .A(arr[1436]), .S(n2928), .Y(n420) );
  MUX2X1 U6387 ( .B(arr[1313]), .A(arr[1354]), .S(n2928), .Y(n419) );
  MUX2X1 U6388 ( .B(n418), .A(n415), .S(n3129), .Y(n422) );
  MUX2X1 U6389 ( .B(n421), .A(n406), .S(n3180), .Y(n455) );
  MUX2X1 U6390 ( .B(arr[1231]), .A(arr[1272]), .S(n2928), .Y(n426) );
  MUX2X1 U6391 ( .B(arr[1149]), .A(arr[1190]), .S(n2928), .Y(n425) );
  MUX2X1 U6392 ( .B(arr[1067]), .A(arr[1108]), .S(n2928), .Y(n429) );
  MUX2X1 U6393 ( .B(arr[985]), .A(arr[1026]), .S(n2928), .Y(n428) );
  MUX2X1 U6394 ( .B(n427), .A(n424), .S(n3129), .Y(n438) );
  MUX2X1 U6395 ( .B(arr[903]), .A(arr[944]), .S(n2929), .Y(n432) );
  MUX2X1 U6396 ( .B(arr[821]), .A(arr[862]), .S(n2929), .Y(n431) );
  MUX2X1 U6397 ( .B(arr[739]), .A(arr[780]), .S(n2929), .Y(n435) );
  MUX2X1 U6398 ( .B(arr[657]), .A(arr[698]), .S(n2929), .Y(n434) );
  MUX2X1 U6399 ( .B(n433), .A(n430), .S(n3129), .Y(n437) );
  MUX2X1 U6400 ( .B(arr[575]), .A(arr[616]), .S(n2929), .Y(n441) );
  MUX2X1 U6401 ( .B(arr[493]), .A(arr[534]), .S(n2929), .Y(n440) );
  MUX2X1 U6402 ( .B(arr[411]), .A(arr[452]), .S(n2929), .Y(n444) );
  MUX2X1 U6403 ( .B(arr[329]), .A(arr[370]), .S(n2929), .Y(n443) );
  MUX2X1 U6404 ( .B(n442), .A(n439), .S(n3129), .Y(n453) );
  MUX2X1 U6405 ( .B(arr[247]), .A(arr[288]), .S(n2929), .Y(n447) );
  MUX2X1 U6406 ( .B(arr[165]), .A(arr[206]), .S(n2929), .Y(n446) );
  MUX2X1 U6407 ( .B(arr[83]), .A(arr[124]), .S(n2929), .Y(n450) );
  MUX2X1 U6408 ( .B(arr[1]), .A(arr[42]), .S(n2929), .Y(n449) );
  MUX2X1 U6409 ( .B(n448), .A(n445), .S(n3129), .Y(n452) );
  MUX2X1 U6410 ( .B(n451), .A(n436), .S(n3180), .Y(n454) );
  MUX2X1 U6411 ( .B(arr[2544]), .A(arr[2585]), .S(n2930), .Y(n458) );
  MUX2X1 U6412 ( .B(arr[2462]), .A(arr[2503]), .S(n2930), .Y(n457) );
  MUX2X1 U6413 ( .B(arr[2380]), .A(arr[2421]), .S(n2930), .Y(n461) );
  MUX2X1 U6414 ( .B(arr[2298]), .A(arr[2339]), .S(n2930), .Y(n460) );
  MUX2X1 U6415 ( .B(n459), .A(n456), .S(n3130), .Y(n470) );
  MUX2X1 U6416 ( .B(arr[2216]), .A(arr[2257]), .S(n2930), .Y(n464) );
  MUX2X1 U6417 ( .B(arr[2134]), .A(arr[2175]), .S(n2930), .Y(n463) );
  MUX2X1 U6418 ( .B(arr[2052]), .A(arr[2093]), .S(n2930), .Y(n467) );
  MUX2X1 U6419 ( .B(arr[1970]), .A(arr[2011]), .S(n2930), .Y(n466) );
  MUX2X1 U6420 ( .B(n465), .A(n462), .S(n3130), .Y(n469) );
  MUX2X1 U6421 ( .B(arr[1888]), .A(arr[1929]), .S(n2930), .Y(n473) );
  MUX2X1 U6422 ( .B(arr[1806]), .A(arr[1847]), .S(n2930), .Y(n472) );
  MUX2X1 U6423 ( .B(arr[1724]), .A(arr[1765]), .S(n2930), .Y(n476) );
  MUX2X1 U6424 ( .B(arr[1642]), .A(arr[1683]), .S(n2930), .Y(n475) );
  MUX2X1 U6425 ( .B(n474), .A(n471), .S(n3130), .Y(n485) );
  MUX2X1 U6426 ( .B(arr[1560]), .A(arr[1601]), .S(n2931), .Y(n479) );
  MUX2X1 U6427 ( .B(arr[1478]), .A(arr[1519]), .S(n2931), .Y(n478) );
  MUX2X1 U6428 ( .B(arr[1396]), .A(arr[1437]), .S(n2931), .Y(n482) );
  MUX2X1 U6429 ( .B(arr[1314]), .A(arr[1355]), .S(n2931), .Y(n481) );
  MUX2X1 U6430 ( .B(n480), .A(n477), .S(n3130), .Y(n484) );
  MUX2X1 U6431 ( .B(n483), .A(n468), .S(n3180), .Y(n517) );
  MUX2X1 U6432 ( .B(arr[1232]), .A(arr[1273]), .S(n2931), .Y(n488) );
  MUX2X1 U6433 ( .B(arr[1150]), .A(arr[1191]), .S(n2931), .Y(n487) );
  MUX2X1 U6434 ( .B(arr[1068]), .A(arr[1109]), .S(n2931), .Y(n491) );
  MUX2X1 U6435 ( .B(arr[986]), .A(arr[1027]), .S(n2931), .Y(n490) );
  MUX2X1 U6436 ( .B(n489), .A(n486), .S(n3130), .Y(n500) );
  MUX2X1 U6437 ( .B(arr[904]), .A(arr[945]), .S(n2931), .Y(n494) );
  MUX2X1 U6438 ( .B(arr[822]), .A(arr[863]), .S(n2931), .Y(n493) );
  MUX2X1 U6439 ( .B(arr[740]), .A(arr[781]), .S(n2931), .Y(n497) );
  MUX2X1 U6440 ( .B(arr[658]), .A(arr[699]), .S(n2931), .Y(n496) );
  MUX2X1 U6441 ( .B(n495), .A(n492), .S(n3130), .Y(n499) );
  MUX2X1 U6442 ( .B(arr[576]), .A(arr[617]), .S(n2932), .Y(n503) );
  MUX2X1 U6443 ( .B(arr[494]), .A(arr[535]), .S(n2932), .Y(n502) );
  MUX2X1 U6444 ( .B(arr[412]), .A(arr[453]), .S(n2932), .Y(n506) );
  MUX2X1 U6445 ( .B(arr[330]), .A(arr[371]), .S(n2932), .Y(n505) );
  MUX2X1 U6446 ( .B(n504), .A(n501), .S(n3130), .Y(n515) );
  MUX2X1 U6447 ( .B(arr[248]), .A(arr[289]), .S(n2932), .Y(n509) );
  MUX2X1 U6448 ( .B(arr[166]), .A(arr[207]), .S(n2932), .Y(n508) );
  MUX2X1 U6449 ( .B(arr[84]), .A(arr[125]), .S(n2932), .Y(n512) );
  MUX2X1 U6450 ( .B(arr[2]), .A(arr[43]), .S(n2932), .Y(n511) );
  MUX2X1 U6451 ( .B(n510), .A(n507), .S(n3130), .Y(n514) );
  MUX2X1 U6452 ( .B(n513), .A(n498), .S(n3180), .Y(n516) );
  MUX2X1 U6453 ( .B(arr[2545]), .A(arr[2586]), .S(n2932), .Y(n520) );
  MUX2X1 U6454 ( .B(arr[2463]), .A(arr[2504]), .S(n2932), .Y(n519) );
  MUX2X1 U6455 ( .B(arr[2381]), .A(arr[2422]), .S(n2932), .Y(n523) );
  MUX2X1 U6456 ( .B(arr[2299]), .A(arr[2340]), .S(n2932), .Y(n522) );
  MUX2X1 U6457 ( .B(n521), .A(n518), .S(n3130), .Y(n532) );
  MUX2X1 U6458 ( .B(arr[2217]), .A(arr[2258]), .S(n2933), .Y(n526) );
  MUX2X1 U6459 ( .B(arr[2135]), .A(arr[2176]), .S(n2933), .Y(n525) );
  MUX2X1 U6460 ( .B(arr[2053]), .A(arr[2094]), .S(n2933), .Y(n529) );
  MUX2X1 U6461 ( .B(arr[1971]), .A(arr[2012]), .S(n2933), .Y(n528) );
  MUX2X1 U6462 ( .B(n527), .A(n524), .S(n3130), .Y(n531) );
  MUX2X1 U6463 ( .B(arr[1889]), .A(arr[1930]), .S(n2933), .Y(n535) );
  MUX2X1 U6464 ( .B(arr[1807]), .A(arr[1848]), .S(n2933), .Y(n534) );
  MUX2X1 U6465 ( .B(arr[1725]), .A(arr[1766]), .S(n2933), .Y(n538) );
  MUX2X1 U6466 ( .B(arr[1643]), .A(arr[1684]), .S(n2933), .Y(n537) );
  MUX2X1 U6467 ( .B(n536), .A(n533), .S(n3130), .Y(n547) );
  MUX2X1 U6468 ( .B(arr[1561]), .A(arr[1602]), .S(n2933), .Y(n541) );
  MUX2X1 U6469 ( .B(arr[1479]), .A(arr[1520]), .S(n2933), .Y(n540) );
  MUX2X1 U6470 ( .B(arr[1397]), .A(arr[1438]), .S(n2933), .Y(n544) );
  MUX2X1 U6471 ( .B(arr[1315]), .A(arr[1356]), .S(n2933), .Y(n543) );
  MUX2X1 U6472 ( .B(n542), .A(n539), .S(n3130), .Y(n546) );
  MUX2X1 U6473 ( .B(n545), .A(n530), .S(n3180), .Y(n579) );
  MUX2X1 U6474 ( .B(arr[1233]), .A(arr[1274]), .S(n2934), .Y(n550) );
  MUX2X1 U6475 ( .B(arr[1151]), .A(arr[1192]), .S(n2934), .Y(n549) );
  MUX2X1 U6476 ( .B(arr[1069]), .A(arr[1110]), .S(n2934), .Y(n553) );
  MUX2X1 U6477 ( .B(arr[987]), .A(arr[1028]), .S(n2934), .Y(n552) );
  MUX2X1 U6478 ( .B(n551), .A(n548), .S(n3131), .Y(n562) );
  MUX2X1 U6479 ( .B(arr[905]), .A(arr[946]), .S(n2934), .Y(n556) );
  MUX2X1 U6480 ( .B(arr[823]), .A(arr[864]), .S(n2934), .Y(n555) );
  MUX2X1 U6481 ( .B(arr[741]), .A(arr[782]), .S(n2934), .Y(n559) );
  MUX2X1 U6482 ( .B(arr[659]), .A(arr[700]), .S(n2934), .Y(n558) );
  MUX2X1 U6483 ( .B(n557), .A(n554), .S(n3131), .Y(n561) );
  MUX2X1 U6484 ( .B(arr[577]), .A(arr[618]), .S(n2934), .Y(n565) );
  MUX2X1 U6485 ( .B(arr[495]), .A(arr[536]), .S(n2934), .Y(n564) );
  MUX2X1 U6486 ( .B(arr[413]), .A(arr[454]), .S(n2934), .Y(n568) );
  MUX2X1 U6487 ( .B(arr[331]), .A(arr[372]), .S(n2934), .Y(n567) );
  MUX2X1 U6488 ( .B(n566), .A(n563), .S(n3131), .Y(n577) );
  MUX2X1 U6489 ( .B(arr[249]), .A(arr[290]), .S(n2935), .Y(n571) );
  MUX2X1 U6490 ( .B(arr[167]), .A(arr[208]), .S(n2935), .Y(n570) );
  MUX2X1 U6491 ( .B(arr[85]), .A(arr[126]), .S(n2935), .Y(n574) );
  MUX2X1 U6492 ( .B(arr[3]), .A(arr[44]), .S(n2935), .Y(n573) );
  MUX2X1 U6493 ( .B(n572), .A(n569), .S(n3131), .Y(n576) );
  MUX2X1 U6494 ( .B(n575), .A(n560), .S(n3180), .Y(n578) );
  MUX2X1 U6495 ( .B(arr[2546]), .A(arr[2587]), .S(n2935), .Y(n582) );
  MUX2X1 U6496 ( .B(arr[2464]), .A(arr[2505]), .S(n2935), .Y(n581) );
  MUX2X1 U6497 ( .B(arr[2382]), .A(arr[2423]), .S(n2935), .Y(n585) );
  MUX2X1 U6498 ( .B(arr[2300]), .A(arr[2341]), .S(n2935), .Y(n584) );
  MUX2X1 U6499 ( .B(n583), .A(n580), .S(n3131), .Y(n594) );
  MUX2X1 U6500 ( .B(arr[2218]), .A(arr[2259]), .S(n2935), .Y(n588) );
  MUX2X1 U6501 ( .B(arr[2136]), .A(arr[2177]), .S(n2935), .Y(n587) );
  MUX2X1 U6502 ( .B(arr[2054]), .A(arr[2095]), .S(n2935), .Y(n591) );
  MUX2X1 U6503 ( .B(arr[1972]), .A(arr[2013]), .S(n2935), .Y(n590) );
  MUX2X1 U6504 ( .B(n589), .A(n586), .S(n3131), .Y(n593) );
  MUX2X1 U6505 ( .B(arr[1890]), .A(arr[1931]), .S(n2936), .Y(n597) );
  MUX2X1 U6506 ( .B(arr[1808]), .A(arr[1849]), .S(n2936), .Y(n596) );
  MUX2X1 U6507 ( .B(arr[1726]), .A(arr[1767]), .S(n2936), .Y(n600) );
  MUX2X1 U6508 ( .B(arr[1644]), .A(arr[1685]), .S(n2936), .Y(n599) );
  MUX2X1 U6509 ( .B(n598), .A(n595), .S(n3131), .Y(n609) );
  MUX2X1 U6510 ( .B(arr[1562]), .A(arr[1603]), .S(n2936), .Y(n603) );
  MUX2X1 U6511 ( .B(arr[1480]), .A(arr[1521]), .S(n2936), .Y(n602) );
  MUX2X1 U6512 ( .B(arr[1398]), .A(arr[1439]), .S(n2936), .Y(n606) );
  MUX2X1 U6513 ( .B(arr[1316]), .A(arr[1357]), .S(n2936), .Y(n605) );
  MUX2X1 U6514 ( .B(n604), .A(n601), .S(n3131), .Y(n608) );
  MUX2X1 U6515 ( .B(n607), .A(n592), .S(n3180), .Y(n641) );
  MUX2X1 U6516 ( .B(arr[1234]), .A(arr[1275]), .S(n2936), .Y(n612) );
  MUX2X1 U6517 ( .B(arr[1152]), .A(arr[1193]), .S(n2936), .Y(n611) );
  MUX2X1 U6518 ( .B(arr[1070]), .A(arr[1111]), .S(n2936), .Y(n615) );
  MUX2X1 U6519 ( .B(arr[988]), .A(arr[1029]), .S(n2936), .Y(n614) );
  MUX2X1 U6520 ( .B(n613), .A(n610), .S(n3131), .Y(n624) );
  MUX2X1 U6521 ( .B(arr[906]), .A(arr[947]), .S(n2937), .Y(n618) );
  MUX2X1 U6522 ( .B(arr[824]), .A(arr[865]), .S(n2937), .Y(n617) );
  MUX2X1 U6523 ( .B(arr[742]), .A(arr[783]), .S(n2937), .Y(n621) );
  MUX2X1 U6524 ( .B(arr[660]), .A(arr[701]), .S(n2937), .Y(n620) );
  MUX2X1 U6525 ( .B(n619), .A(n616), .S(n3131), .Y(n623) );
  MUX2X1 U6526 ( .B(arr[578]), .A(arr[619]), .S(n2937), .Y(n627) );
  MUX2X1 U6527 ( .B(arr[496]), .A(arr[537]), .S(n2937), .Y(n626) );
  MUX2X1 U6528 ( .B(arr[414]), .A(arr[455]), .S(n2937), .Y(n630) );
  MUX2X1 U6529 ( .B(arr[332]), .A(arr[373]), .S(n2937), .Y(n629) );
  MUX2X1 U6530 ( .B(n628), .A(n625), .S(n3131), .Y(n639) );
  MUX2X1 U6531 ( .B(arr[250]), .A(arr[291]), .S(n2937), .Y(n633) );
  MUX2X1 U6532 ( .B(arr[168]), .A(arr[209]), .S(n2937), .Y(n632) );
  MUX2X1 U6533 ( .B(arr[86]), .A(arr[127]), .S(n2937), .Y(n636) );
  MUX2X1 U6534 ( .B(arr[4]), .A(arr[45]), .S(n2937), .Y(n635) );
  MUX2X1 U6535 ( .B(n634), .A(n631), .S(n3131), .Y(n638) );
  MUX2X1 U6536 ( .B(n637), .A(n622), .S(n3180), .Y(n640) );
  MUX2X1 U6537 ( .B(arr[2547]), .A(arr[2588]), .S(n2938), .Y(n644) );
  MUX2X1 U6538 ( .B(arr[2465]), .A(arr[2506]), .S(n2938), .Y(n643) );
  MUX2X1 U6539 ( .B(arr[2383]), .A(arr[2424]), .S(n2938), .Y(n647) );
  MUX2X1 U6540 ( .B(arr[2301]), .A(arr[2342]), .S(n2938), .Y(n646) );
  MUX2X1 U6541 ( .B(n645), .A(n642), .S(n3132), .Y(n656) );
  MUX2X1 U6542 ( .B(arr[2219]), .A(arr[2260]), .S(n2938), .Y(n650) );
  MUX2X1 U6543 ( .B(arr[2137]), .A(arr[2178]), .S(n2938), .Y(n649) );
  MUX2X1 U6544 ( .B(arr[2055]), .A(arr[2096]), .S(n2938), .Y(n653) );
  MUX2X1 U6545 ( .B(arr[1973]), .A(arr[2014]), .S(n2938), .Y(n652) );
  MUX2X1 U6546 ( .B(n651), .A(n648), .S(n3132), .Y(n655) );
  MUX2X1 U6547 ( .B(arr[1891]), .A(arr[1932]), .S(n2938), .Y(n659) );
  MUX2X1 U6548 ( .B(arr[1809]), .A(arr[1850]), .S(n2938), .Y(n658) );
  MUX2X1 U6549 ( .B(arr[1727]), .A(arr[1768]), .S(n2938), .Y(n662) );
  MUX2X1 U6550 ( .B(arr[1645]), .A(arr[1686]), .S(n2938), .Y(n661) );
  MUX2X1 U6551 ( .B(n660), .A(n657), .S(n3132), .Y(n671) );
  MUX2X1 U6552 ( .B(arr[1563]), .A(arr[1604]), .S(n2939), .Y(n665) );
  MUX2X1 U6553 ( .B(arr[1481]), .A(arr[1522]), .S(n2939), .Y(n664) );
  MUX2X1 U6554 ( .B(arr[1399]), .A(arr[1440]), .S(n2939), .Y(n668) );
  MUX2X1 U6555 ( .B(arr[1317]), .A(arr[1358]), .S(n2939), .Y(n667) );
  MUX2X1 U6556 ( .B(n666), .A(n663), .S(n3132), .Y(n670) );
  MUX2X1 U6557 ( .B(n669), .A(n654), .S(n3181), .Y(n703) );
  MUX2X1 U6558 ( .B(arr[1235]), .A(arr[1276]), .S(n2939), .Y(n674) );
  MUX2X1 U6559 ( .B(arr[1153]), .A(arr[1194]), .S(n2939), .Y(n673) );
  MUX2X1 U6560 ( .B(arr[1071]), .A(arr[1112]), .S(n2939), .Y(n677) );
  MUX2X1 U6561 ( .B(arr[989]), .A(arr[1030]), .S(n2939), .Y(n676) );
  MUX2X1 U6562 ( .B(n675), .A(n672), .S(n3132), .Y(n686) );
  MUX2X1 U6563 ( .B(arr[907]), .A(arr[948]), .S(n2939), .Y(n680) );
  MUX2X1 U6564 ( .B(arr[825]), .A(arr[866]), .S(n2939), .Y(n679) );
  MUX2X1 U6565 ( .B(arr[743]), .A(arr[784]), .S(n2939), .Y(n683) );
  MUX2X1 U6566 ( .B(arr[661]), .A(arr[702]), .S(n2939), .Y(n682) );
  MUX2X1 U6567 ( .B(n681), .A(n678), .S(n3132), .Y(n685) );
  MUX2X1 U6568 ( .B(arr[579]), .A(arr[620]), .S(n2940), .Y(n689) );
  MUX2X1 U6569 ( .B(arr[497]), .A(arr[538]), .S(n2940), .Y(n688) );
  MUX2X1 U6570 ( .B(arr[415]), .A(arr[456]), .S(n2940), .Y(n692) );
  MUX2X1 U6571 ( .B(arr[333]), .A(arr[374]), .S(n2940), .Y(n691) );
  MUX2X1 U6572 ( .B(n690), .A(n687), .S(n3132), .Y(n701) );
  MUX2X1 U6573 ( .B(arr[251]), .A(arr[292]), .S(n2940), .Y(n695) );
  MUX2X1 U6574 ( .B(arr[169]), .A(arr[210]), .S(n2940), .Y(n694) );
  MUX2X1 U6575 ( .B(arr[87]), .A(arr[128]), .S(n2940), .Y(n698) );
  MUX2X1 U6576 ( .B(arr[5]), .A(arr[46]), .S(n2940), .Y(n697) );
  MUX2X1 U6577 ( .B(n696), .A(n693), .S(n3132), .Y(n700) );
  MUX2X1 U6578 ( .B(n699), .A(n684), .S(n3181), .Y(n702) );
  MUX2X1 U6579 ( .B(arr[2548]), .A(arr[2589]), .S(n2940), .Y(n706) );
  MUX2X1 U6580 ( .B(arr[2466]), .A(arr[2507]), .S(n2940), .Y(n705) );
  MUX2X1 U6581 ( .B(arr[2384]), .A(arr[2425]), .S(n2940), .Y(n709) );
  MUX2X1 U6582 ( .B(arr[2302]), .A(arr[2343]), .S(n2940), .Y(n708) );
  MUX2X1 U6583 ( .B(n707), .A(n704), .S(n3132), .Y(n718) );
  MUX2X1 U6584 ( .B(arr[2220]), .A(arr[2261]), .S(n2941), .Y(n712) );
  MUX2X1 U6585 ( .B(arr[2138]), .A(arr[2179]), .S(n2941), .Y(n711) );
  MUX2X1 U6586 ( .B(arr[2056]), .A(arr[2097]), .S(n2941), .Y(n715) );
  MUX2X1 U6587 ( .B(arr[1974]), .A(arr[2015]), .S(n2941), .Y(n714) );
  MUX2X1 U6588 ( .B(n713), .A(n710), .S(n3132), .Y(n717) );
  MUX2X1 U6589 ( .B(arr[1892]), .A(arr[1933]), .S(n2941), .Y(n721) );
  MUX2X1 U6590 ( .B(arr[1810]), .A(arr[1851]), .S(n2941), .Y(n720) );
  MUX2X1 U6591 ( .B(arr[1728]), .A(arr[1769]), .S(n2941), .Y(n724) );
  MUX2X1 U6592 ( .B(arr[1646]), .A(arr[1687]), .S(n2941), .Y(n723) );
  MUX2X1 U6593 ( .B(n722), .A(n719), .S(n3132), .Y(n733) );
  MUX2X1 U6594 ( .B(arr[1564]), .A(arr[1605]), .S(n2941), .Y(n727) );
  MUX2X1 U6595 ( .B(arr[1482]), .A(arr[1523]), .S(n2941), .Y(n726) );
  MUX2X1 U6596 ( .B(arr[1400]), .A(arr[1441]), .S(n2941), .Y(n730) );
  MUX2X1 U6597 ( .B(arr[1318]), .A(arr[1359]), .S(n2941), .Y(n729) );
  MUX2X1 U6598 ( .B(n728), .A(n725), .S(n3132), .Y(n732) );
  MUX2X1 U6599 ( .B(n731), .A(n716), .S(n3181), .Y(n765) );
  MUX2X1 U6600 ( .B(arr[1236]), .A(arr[1277]), .S(n2942), .Y(n736) );
  MUX2X1 U6601 ( .B(arr[1154]), .A(arr[1195]), .S(n2942), .Y(n735) );
  MUX2X1 U6602 ( .B(arr[1072]), .A(arr[1113]), .S(n2942), .Y(n739) );
  MUX2X1 U6603 ( .B(arr[990]), .A(arr[1031]), .S(n2942), .Y(n738) );
  MUX2X1 U6604 ( .B(n737), .A(n734), .S(n3133), .Y(n748) );
  MUX2X1 U6605 ( .B(arr[908]), .A(arr[949]), .S(n2942), .Y(n742) );
  MUX2X1 U6606 ( .B(arr[826]), .A(arr[867]), .S(n2942), .Y(n741) );
  MUX2X1 U6607 ( .B(arr[744]), .A(arr[785]), .S(n2942), .Y(n745) );
  MUX2X1 U6608 ( .B(arr[662]), .A(arr[703]), .S(n2942), .Y(n744) );
  MUX2X1 U6609 ( .B(n743), .A(n740), .S(n3133), .Y(n747) );
  MUX2X1 U6610 ( .B(arr[580]), .A(arr[621]), .S(n2942), .Y(n751) );
  MUX2X1 U6611 ( .B(arr[498]), .A(arr[539]), .S(n2942), .Y(n750) );
  MUX2X1 U6612 ( .B(arr[416]), .A(arr[457]), .S(n2942), .Y(n754) );
  MUX2X1 U6613 ( .B(arr[334]), .A(arr[375]), .S(n2942), .Y(n753) );
  MUX2X1 U6614 ( .B(n752), .A(n749), .S(n3133), .Y(n763) );
  MUX2X1 U6615 ( .B(arr[252]), .A(arr[293]), .S(n2943), .Y(n757) );
  MUX2X1 U6616 ( .B(arr[170]), .A(arr[211]), .S(n2943), .Y(n756) );
  MUX2X1 U6617 ( .B(arr[88]), .A(arr[129]), .S(n2943), .Y(n760) );
  MUX2X1 U6618 ( .B(arr[6]), .A(arr[47]), .S(n2943), .Y(n759) );
  MUX2X1 U6619 ( .B(n758), .A(n755), .S(n3133), .Y(n762) );
  MUX2X1 U6620 ( .B(n761), .A(n746), .S(n3181), .Y(n764) );
  MUX2X1 U6621 ( .B(arr[2549]), .A(arr[2590]), .S(n2943), .Y(n768) );
  MUX2X1 U6622 ( .B(arr[2467]), .A(arr[2508]), .S(n2943), .Y(n767) );
  MUX2X1 U6623 ( .B(arr[2385]), .A(arr[2426]), .S(n2943), .Y(n771) );
  MUX2X1 U6624 ( .B(arr[2303]), .A(arr[2344]), .S(n2943), .Y(n770) );
  MUX2X1 U6625 ( .B(n769), .A(n766), .S(n3133), .Y(n780) );
  MUX2X1 U6626 ( .B(arr[2221]), .A(arr[2262]), .S(n2943), .Y(n774) );
  MUX2X1 U6627 ( .B(arr[2139]), .A(arr[2180]), .S(n2943), .Y(n773) );
  MUX2X1 U6628 ( .B(arr[2057]), .A(arr[2098]), .S(n2943), .Y(n777) );
  MUX2X1 U6629 ( .B(arr[1975]), .A(arr[2016]), .S(n2943), .Y(n776) );
  MUX2X1 U6630 ( .B(n775), .A(n772), .S(n3133), .Y(n779) );
  MUX2X1 U6631 ( .B(arr[1893]), .A(arr[1934]), .S(n2944), .Y(n783) );
  MUX2X1 U6632 ( .B(arr[1811]), .A(arr[1852]), .S(n2944), .Y(n782) );
  MUX2X1 U6633 ( .B(arr[1729]), .A(arr[1770]), .S(n2944), .Y(n786) );
  MUX2X1 U6634 ( .B(arr[1647]), .A(arr[1688]), .S(n2944), .Y(n785) );
  MUX2X1 U6635 ( .B(n784), .A(n781), .S(n3133), .Y(n795) );
  MUX2X1 U6636 ( .B(arr[1565]), .A(arr[1606]), .S(n2944), .Y(n789) );
  MUX2X1 U6637 ( .B(arr[1483]), .A(arr[1524]), .S(n2944), .Y(n788) );
  MUX2X1 U6638 ( .B(arr[1401]), .A(arr[1442]), .S(n2944), .Y(n792) );
  MUX2X1 U6639 ( .B(arr[1319]), .A(arr[1360]), .S(n2944), .Y(n791) );
  MUX2X1 U6640 ( .B(n790), .A(n787), .S(n3133), .Y(n794) );
  MUX2X1 U6641 ( .B(n793), .A(n778), .S(n3181), .Y(n827) );
  MUX2X1 U6642 ( .B(arr[1237]), .A(arr[1278]), .S(n2944), .Y(n798) );
  MUX2X1 U6643 ( .B(arr[1155]), .A(arr[1196]), .S(n2944), .Y(n797) );
  MUX2X1 U6644 ( .B(arr[1073]), .A(arr[1114]), .S(n2944), .Y(n801) );
  MUX2X1 U6645 ( .B(arr[991]), .A(arr[1032]), .S(n2944), .Y(n800) );
  MUX2X1 U6646 ( .B(n799), .A(n796), .S(n3133), .Y(n810) );
  MUX2X1 U6647 ( .B(arr[909]), .A(arr[950]), .S(n2945), .Y(n804) );
  MUX2X1 U6648 ( .B(arr[827]), .A(arr[868]), .S(n2945), .Y(n803) );
  MUX2X1 U6649 ( .B(arr[745]), .A(arr[786]), .S(n2945), .Y(n807) );
  MUX2X1 U6650 ( .B(arr[663]), .A(arr[704]), .S(n2945), .Y(n806) );
  MUX2X1 U6651 ( .B(n805), .A(n802), .S(n3133), .Y(n809) );
  MUX2X1 U6652 ( .B(arr[581]), .A(arr[622]), .S(n2945), .Y(n813) );
  MUX2X1 U6653 ( .B(arr[499]), .A(arr[540]), .S(n2945), .Y(n812) );
  MUX2X1 U6654 ( .B(arr[417]), .A(arr[458]), .S(n2945), .Y(n816) );
  MUX2X1 U6655 ( .B(arr[335]), .A(arr[376]), .S(n2945), .Y(n815) );
  MUX2X1 U6656 ( .B(n814), .A(n811), .S(n3133), .Y(n825) );
  MUX2X1 U6657 ( .B(arr[253]), .A(arr[294]), .S(n2945), .Y(n819) );
  MUX2X1 U6658 ( .B(arr[171]), .A(arr[212]), .S(n2945), .Y(n818) );
  MUX2X1 U6659 ( .B(arr[89]), .A(arr[130]), .S(n2945), .Y(n822) );
  MUX2X1 U6660 ( .B(arr[7]), .A(arr[48]), .S(n2945), .Y(n821) );
  MUX2X1 U6661 ( .B(n820), .A(n817), .S(n3133), .Y(n824) );
  MUX2X1 U6662 ( .B(n823), .A(n808), .S(n3181), .Y(n826) );
  MUX2X1 U6663 ( .B(arr[2550]), .A(arr[2591]), .S(n2946), .Y(n830) );
  MUX2X1 U6664 ( .B(arr[2468]), .A(arr[2509]), .S(n2946), .Y(n829) );
  MUX2X1 U6665 ( .B(arr[2386]), .A(arr[2427]), .S(n2946), .Y(n833) );
  MUX2X1 U6666 ( .B(arr[2304]), .A(arr[2345]), .S(n2946), .Y(n832) );
  MUX2X1 U6667 ( .B(n831), .A(n828), .S(n3134), .Y(n842) );
  MUX2X1 U6668 ( .B(arr[2222]), .A(arr[2263]), .S(n2946), .Y(n836) );
  MUX2X1 U6669 ( .B(arr[2140]), .A(arr[2181]), .S(n2946), .Y(n835) );
  MUX2X1 U6670 ( .B(arr[2058]), .A(arr[2099]), .S(n2946), .Y(n839) );
  MUX2X1 U6671 ( .B(arr[1976]), .A(arr[2017]), .S(n2946), .Y(n838) );
  MUX2X1 U6672 ( .B(n837), .A(n834), .S(n3134), .Y(n841) );
  MUX2X1 U6673 ( .B(arr[1894]), .A(arr[1935]), .S(n2946), .Y(n845) );
  MUX2X1 U6674 ( .B(arr[1812]), .A(arr[1853]), .S(n2946), .Y(n844) );
  MUX2X1 U6675 ( .B(arr[1730]), .A(arr[1771]), .S(n2946), .Y(n848) );
  MUX2X1 U6676 ( .B(arr[1648]), .A(arr[1689]), .S(n2946), .Y(n847) );
  MUX2X1 U6677 ( .B(n846), .A(n843), .S(n3134), .Y(n857) );
  MUX2X1 U6678 ( .B(arr[1566]), .A(arr[1607]), .S(n2947), .Y(n851) );
  MUX2X1 U6679 ( .B(arr[1484]), .A(arr[1525]), .S(n2947), .Y(n850) );
  MUX2X1 U6680 ( .B(arr[1402]), .A(arr[1443]), .S(n2947), .Y(n854) );
  MUX2X1 U6681 ( .B(arr[1320]), .A(arr[1361]), .S(n2947), .Y(n853) );
  MUX2X1 U6682 ( .B(n852), .A(n849), .S(n3134), .Y(n856) );
  MUX2X1 U6683 ( .B(n855), .A(n840), .S(n3181), .Y(n889) );
  MUX2X1 U6684 ( .B(arr[1238]), .A(arr[1279]), .S(n2947), .Y(n860) );
  MUX2X1 U6685 ( .B(arr[1156]), .A(arr[1197]), .S(n2947), .Y(n859) );
  MUX2X1 U6686 ( .B(arr[1074]), .A(arr[1115]), .S(n2947), .Y(n863) );
  MUX2X1 U6687 ( .B(arr[992]), .A(arr[1033]), .S(n2947), .Y(n862) );
  MUX2X1 U6688 ( .B(n861), .A(n858), .S(n3134), .Y(n872) );
  MUX2X1 U6689 ( .B(arr[910]), .A(arr[951]), .S(n2947), .Y(n866) );
  MUX2X1 U6690 ( .B(arr[828]), .A(arr[869]), .S(n2947), .Y(n865) );
  MUX2X1 U6691 ( .B(arr[746]), .A(arr[787]), .S(n2947), .Y(n869) );
  MUX2X1 U6692 ( .B(arr[664]), .A(arr[705]), .S(n2947), .Y(n868) );
  MUX2X1 U6693 ( .B(n867), .A(n864), .S(n3134), .Y(n871) );
  MUX2X1 U6694 ( .B(arr[582]), .A(arr[623]), .S(n2948), .Y(n875) );
  MUX2X1 U6695 ( .B(arr[500]), .A(arr[541]), .S(n2948), .Y(n874) );
  MUX2X1 U6696 ( .B(arr[418]), .A(arr[459]), .S(n2948), .Y(n878) );
  MUX2X1 U6697 ( .B(arr[336]), .A(arr[377]), .S(n2948), .Y(n877) );
  MUX2X1 U6698 ( .B(n876), .A(n873), .S(n3134), .Y(n887) );
  MUX2X1 U6699 ( .B(arr[254]), .A(arr[295]), .S(n2948), .Y(n881) );
  MUX2X1 U6700 ( .B(arr[172]), .A(arr[213]), .S(n2948), .Y(n880) );
  MUX2X1 U6701 ( .B(arr[90]), .A(arr[131]), .S(n2948), .Y(n884) );
  MUX2X1 U6702 ( .B(arr[8]), .A(arr[49]), .S(n2948), .Y(n883) );
  MUX2X1 U6703 ( .B(n882), .A(n879), .S(n3134), .Y(n886) );
  MUX2X1 U6704 ( .B(n885), .A(n870), .S(n3181), .Y(n888) );
  MUX2X1 U6705 ( .B(arr[2551]), .A(arr[2592]), .S(n2948), .Y(n892) );
  MUX2X1 U6706 ( .B(arr[2469]), .A(arr[2510]), .S(n2948), .Y(n891) );
  MUX2X1 U6707 ( .B(arr[2387]), .A(arr[2428]), .S(n2948), .Y(n895) );
  MUX2X1 U6708 ( .B(arr[2305]), .A(arr[2346]), .S(n2948), .Y(n894) );
  MUX2X1 U6709 ( .B(n893), .A(n890), .S(n3134), .Y(n904) );
  MUX2X1 U6710 ( .B(arr[2223]), .A(arr[2264]), .S(n2949), .Y(n898) );
  MUX2X1 U6711 ( .B(arr[2141]), .A(arr[2182]), .S(n2949), .Y(n897) );
  MUX2X1 U6712 ( .B(arr[2059]), .A(arr[2100]), .S(n2949), .Y(n901) );
  MUX2X1 U6713 ( .B(arr[1977]), .A(arr[2018]), .S(n2949), .Y(n900) );
  MUX2X1 U6714 ( .B(n899), .A(n896), .S(n3134), .Y(n903) );
  MUX2X1 U6715 ( .B(arr[1895]), .A(arr[1936]), .S(n2949), .Y(n907) );
  MUX2X1 U6716 ( .B(arr[1813]), .A(arr[1854]), .S(n2949), .Y(n906) );
  MUX2X1 U6717 ( .B(arr[1731]), .A(arr[1772]), .S(n2949), .Y(n910) );
  MUX2X1 U6718 ( .B(arr[1649]), .A(arr[1690]), .S(n2949), .Y(n909) );
  MUX2X1 U6719 ( .B(n908), .A(n905), .S(n3134), .Y(n919) );
  MUX2X1 U6720 ( .B(arr[1567]), .A(arr[1608]), .S(n2949), .Y(n913) );
  MUX2X1 U6721 ( .B(arr[1485]), .A(arr[1526]), .S(n2949), .Y(n912) );
  MUX2X1 U6722 ( .B(arr[1403]), .A(arr[1444]), .S(n2949), .Y(n916) );
  MUX2X1 U6723 ( .B(arr[1321]), .A(arr[1362]), .S(n2949), .Y(n915) );
  MUX2X1 U6724 ( .B(n914), .A(n911), .S(n3134), .Y(n918) );
  MUX2X1 U6725 ( .B(n917), .A(n902), .S(n3181), .Y(n951) );
  MUX2X1 U6726 ( .B(arr[1239]), .A(arr[1280]), .S(n2950), .Y(n922) );
  MUX2X1 U6727 ( .B(arr[1157]), .A(arr[1198]), .S(n2950), .Y(n921) );
  MUX2X1 U6728 ( .B(arr[1075]), .A(arr[1116]), .S(n2950), .Y(n925) );
  MUX2X1 U6729 ( .B(arr[993]), .A(arr[1034]), .S(n2950), .Y(n924) );
  MUX2X1 U6730 ( .B(n923), .A(n920), .S(n3135), .Y(n934) );
  MUX2X1 U6731 ( .B(arr[911]), .A(arr[952]), .S(n2950), .Y(n928) );
  MUX2X1 U6732 ( .B(arr[829]), .A(arr[870]), .S(n2950), .Y(n927) );
  MUX2X1 U6733 ( .B(arr[747]), .A(arr[788]), .S(n2950), .Y(n931) );
  MUX2X1 U6734 ( .B(arr[665]), .A(arr[706]), .S(n2950), .Y(n930) );
  MUX2X1 U6735 ( .B(n929), .A(n926), .S(n3135), .Y(n933) );
  MUX2X1 U6736 ( .B(arr[583]), .A(arr[624]), .S(n2950), .Y(n937) );
  MUX2X1 U6737 ( .B(arr[501]), .A(arr[542]), .S(n2950), .Y(n936) );
  MUX2X1 U6738 ( .B(arr[419]), .A(arr[460]), .S(n2950), .Y(n940) );
  MUX2X1 U6739 ( .B(arr[337]), .A(arr[378]), .S(n2950), .Y(n939) );
  MUX2X1 U6740 ( .B(n938), .A(n935), .S(n3135), .Y(n949) );
  MUX2X1 U6741 ( .B(arr[255]), .A(arr[296]), .S(n2951), .Y(n943) );
  MUX2X1 U6742 ( .B(arr[173]), .A(arr[214]), .S(n2951), .Y(n942) );
  MUX2X1 U6743 ( .B(arr[91]), .A(arr[132]), .S(n2951), .Y(n946) );
  MUX2X1 U6744 ( .B(arr[9]), .A(arr[50]), .S(n2951), .Y(n945) );
  MUX2X1 U6745 ( .B(n944), .A(n941), .S(n3135), .Y(n948) );
  MUX2X1 U6746 ( .B(n947), .A(n932), .S(n3181), .Y(n950) );
  MUX2X1 U6747 ( .B(arr[2552]), .A(arr[2593]), .S(n2951), .Y(n954) );
  MUX2X1 U6748 ( .B(arr[2470]), .A(arr[2511]), .S(n2951), .Y(n953) );
  MUX2X1 U6749 ( .B(arr[2388]), .A(arr[2429]), .S(n2951), .Y(n957) );
  MUX2X1 U6750 ( .B(arr[2306]), .A(arr[2347]), .S(n2951), .Y(n956) );
  MUX2X1 U6751 ( .B(n955), .A(n952), .S(n3135), .Y(n966) );
  MUX2X1 U6752 ( .B(arr[2224]), .A(arr[2265]), .S(n2951), .Y(n960) );
  MUX2X1 U6753 ( .B(arr[2142]), .A(arr[2183]), .S(n2951), .Y(n959) );
  MUX2X1 U6754 ( .B(arr[2060]), .A(arr[2101]), .S(n2951), .Y(n963) );
  MUX2X1 U6755 ( .B(arr[1978]), .A(arr[2019]), .S(n2951), .Y(n962) );
  MUX2X1 U6756 ( .B(n961), .A(n958), .S(n3135), .Y(n965) );
  MUX2X1 U6757 ( .B(arr[1896]), .A(arr[1937]), .S(n2952), .Y(n969) );
  MUX2X1 U6758 ( .B(arr[1814]), .A(arr[1855]), .S(n2952), .Y(n968) );
  MUX2X1 U6759 ( .B(arr[1732]), .A(arr[1773]), .S(n2952), .Y(n972) );
  MUX2X1 U6760 ( .B(arr[1650]), .A(arr[1691]), .S(n2952), .Y(n971) );
  MUX2X1 U6761 ( .B(n970), .A(n967), .S(n3135), .Y(n981) );
  MUX2X1 U6762 ( .B(arr[1568]), .A(arr[1609]), .S(n2952), .Y(n975) );
  MUX2X1 U6763 ( .B(arr[1486]), .A(arr[1527]), .S(n2952), .Y(n974) );
  MUX2X1 U6764 ( .B(arr[1404]), .A(arr[1445]), .S(n2952), .Y(n978) );
  MUX2X1 U6765 ( .B(arr[1322]), .A(arr[1363]), .S(n2952), .Y(n977) );
  MUX2X1 U6766 ( .B(n976), .A(n973), .S(n3135), .Y(n980) );
  MUX2X1 U6767 ( .B(n979), .A(n964), .S(n3181), .Y(n1013) );
  MUX2X1 U6768 ( .B(arr[1240]), .A(arr[1281]), .S(n2952), .Y(n984) );
  MUX2X1 U6769 ( .B(arr[1158]), .A(arr[1199]), .S(n2952), .Y(n983) );
  MUX2X1 U6770 ( .B(arr[1076]), .A(arr[1117]), .S(n2952), .Y(n987) );
  MUX2X1 U6771 ( .B(arr[994]), .A(arr[1035]), .S(n2952), .Y(n986) );
  MUX2X1 U6772 ( .B(n985), .A(n982), .S(n3135), .Y(n996) );
  MUX2X1 U6773 ( .B(arr[912]), .A(arr[953]), .S(n2953), .Y(n990) );
  MUX2X1 U6774 ( .B(arr[830]), .A(arr[871]), .S(n2953), .Y(n989) );
  MUX2X1 U6775 ( .B(arr[748]), .A(arr[789]), .S(n2953), .Y(n993) );
  MUX2X1 U6776 ( .B(arr[666]), .A(arr[707]), .S(n2953), .Y(n992) );
  MUX2X1 U6777 ( .B(n991), .A(n988), .S(n3135), .Y(n995) );
  MUX2X1 U6778 ( .B(arr[584]), .A(arr[625]), .S(n2953), .Y(n999) );
  MUX2X1 U6779 ( .B(arr[502]), .A(arr[543]), .S(n2953), .Y(n998) );
  MUX2X1 U6780 ( .B(arr[420]), .A(arr[461]), .S(n2953), .Y(n1002) );
  MUX2X1 U6781 ( .B(arr[338]), .A(arr[379]), .S(n2953), .Y(n1001) );
  MUX2X1 U6782 ( .B(n1000), .A(n997), .S(n3135), .Y(n1011) );
  MUX2X1 U6783 ( .B(arr[256]), .A(arr[297]), .S(n2953), .Y(n1005) );
  MUX2X1 U6784 ( .B(arr[174]), .A(arr[215]), .S(n2953), .Y(n1004) );
  MUX2X1 U6785 ( .B(arr[92]), .A(arr[133]), .S(n2953), .Y(n1008) );
  MUX2X1 U6786 ( .B(arr[10]), .A(arr[51]), .S(n2953), .Y(n1007) );
  MUX2X1 U6787 ( .B(n1006), .A(n1003), .S(n3135), .Y(n1010) );
  MUX2X1 U6788 ( .B(n1009), .A(n994), .S(n3181), .Y(n1012) );
  MUX2X1 U6789 ( .B(arr[2553]), .A(arr[2594]), .S(n2954), .Y(n1016) );
  MUX2X1 U6790 ( .B(arr[2471]), .A(arr[2512]), .S(n2954), .Y(n1015) );
  MUX2X1 U6791 ( .B(arr[2389]), .A(arr[2430]), .S(n2954), .Y(n1019) );
  MUX2X1 U6792 ( .B(arr[2307]), .A(arr[2348]), .S(n2954), .Y(n1018) );
  MUX2X1 U6793 ( .B(n1017), .A(n1014), .S(n3136), .Y(n1028) );
  MUX2X1 U6794 ( .B(arr[2225]), .A(arr[2266]), .S(n2954), .Y(n1022) );
  MUX2X1 U6795 ( .B(arr[2143]), .A(arr[2184]), .S(n2954), .Y(n1021) );
  MUX2X1 U6796 ( .B(arr[2061]), .A(arr[2102]), .S(n2954), .Y(n1025) );
  MUX2X1 U6797 ( .B(arr[1979]), .A(arr[2020]), .S(n2954), .Y(n1024) );
  MUX2X1 U6798 ( .B(n1023), .A(n1020), .S(n3136), .Y(n1027) );
  MUX2X1 U6799 ( .B(arr[1897]), .A(arr[1938]), .S(n2954), .Y(n1031) );
  MUX2X1 U6800 ( .B(arr[1815]), .A(arr[1856]), .S(n2954), .Y(n1030) );
  MUX2X1 U6801 ( .B(arr[1733]), .A(arr[1774]), .S(n2954), .Y(n1034) );
  MUX2X1 U6802 ( .B(arr[1651]), .A(arr[1692]), .S(n2954), .Y(n1033) );
  MUX2X1 U6803 ( .B(n1032), .A(n1029), .S(n3136), .Y(n1043) );
  MUX2X1 U6804 ( .B(arr[1569]), .A(arr[1610]), .S(n2955), .Y(n1037) );
  MUX2X1 U6805 ( .B(arr[1487]), .A(arr[1528]), .S(n2955), .Y(n1036) );
  MUX2X1 U6806 ( .B(arr[1405]), .A(arr[1446]), .S(n2955), .Y(n1040) );
  MUX2X1 U6807 ( .B(arr[1323]), .A(arr[1364]), .S(n2955), .Y(n1039) );
  MUX2X1 U6808 ( .B(n1038), .A(n1035), .S(n3136), .Y(n1042) );
  MUX2X1 U6809 ( .B(n1041), .A(n1026), .S(n3182), .Y(n1075) );
  MUX2X1 U6810 ( .B(arr[1241]), .A(arr[1282]), .S(n2955), .Y(n1046) );
  MUX2X1 U6811 ( .B(arr[1159]), .A(arr[1200]), .S(n2955), .Y(n1045) );
  MUX2X1 U6812 ( .B(arr[1077]), .A(arr[1118]), .S(n2955), .Y(n1049) );
  MUX2X1 U6813 ( .B(arr[995]), .A(arr[1036]), .S(n2955), .Y(n1048) );
  MUX2X1 U6814 ( .B(n1047), .A(n1044), .S(n3136), .Y(n1058) );
  MUX2X1 U6815 ( .B(arr[913]), .A(arr[954]), .S(n2955), .Y(n1052) );
  MUX2X1 U6816 ( .B(arr[831]), .A(arr[872]), .S(n2955), .Y(n1051) );
  MUX2X1 U6817 ( .B(arr[749]), .A(arr[790]), .S(n2955), .Y(n1055) );
  MUX2X1 U6818 ( .B(arr[667]), .A(arr[708]), .S(n2955), .Y(n1054) );
  MUX2X1 U6819 ( .B(n1053), .A(n1050), .S(n3136), .Y(n1057) );
  MUX2X1 U6820 ( .B(arr[585]), .A(arr[626]), .S(n2956), .Y(n1061) );
  MUX2X1 U6821 ( .B(arr[503]), .A(arr[544]), .S(n2956), .Y(n1060) );
  MUX2X1 U6822 ( .B(arr[421]), .A(arr[462]), .S(n2956), .Y(n1064) );
  MUX2X1 U6823 ( .B(arr[339]), .A(arr[380]), .S(n2956), .Y(n1063) );
  MUX2X1 U6824 ( .B(n1062), .A(n1059), .S(n3136), .Y(n1073) );
  MUX2X1 U6825 ( .B(arr[257]), .A(arr[298]), .S(n2956), .Y(n1067) );
  MUX2X1 U6826 ( .B(arr[175]), .A(arr[216]), .S(n2956), .Y(n1066) );
  MUX2X1 U6827 ( .B(arr[93]), .A(arr[134]), .S(n2956), .Y(n1070) );
  MUX2X1 U6828 ( .B(arr[11]), .A(arr[52]), .S(n2956), .Y(n1069) );
  MUX2X1 U6829 ( .B(n1068), .A(n1065), .S(n3136), .Y(n1072) );
  MUX2X1 U6830 ( .B(n1071), .A(n1056), .S(n3182), .Y(n1074) );
  MUX2X1 U6831 ( .B(arr[2554]), .A(arr[2595]), .S(n2956), .Y(n1078) );
  MUX2X1 U6832 ( .B(arr[2472]), .A(arr[2513]), .S(n2956), .Y(n1077) );
  MUX2X1 U6833 ( .B(arr[2390]), .A(arr[2431]), .S(n2956), .Y(n1081) );
  MUX2X1 U6834 ( .B(arr[2308]), .A(arr[2349]), .S(n2956), .Y(n1080) );
  MUX2X1 U6835 ( .B(n1079), .A(n1076), .S(n3136), .Y(n1090) );
  MUX2X1 U6836 ( .B(arr[2226]), .A(arr[2267]), .S(n2957), .Y(n1084) );
  MUX2X1 U6837 ( .B(arr[2144]), .A(arr[2185]), .S(n2957), .Y(n1083) );
  MUX2X1 U6838 ( .B(arr[2062]), .A(arr[2103]), .S(n2957), .Y(n1087) );
  MUX2X1 U6839 ( .B(arr[1980]), .A(arr[2021]), .S(n2957), .Y(n1086) );
  MUX2X1 U6840 ( .B(n1085), .A(n1082), .S(n3136), .Y(n1089) );
  MUX2X1 U6841 ( .B(arr[1898]), .A(arr[1939]), .S(n2957), .Y(n1093) );
  MUX2X1 U6842 ( .B(arr[1816]), .A(arr[1857]), .S(n2957), .Y(n1092) );
  MUX2X1 U6843 ( .B(arr[1734]), .A(arr[1775]), .S(n2957), .Y(n1096) );
  MUX2X1 U6844 ( .B(arr[1652]), .A(arr[1693]), .S(n2957), .Y(n1095) );
  MUX2X1 U6845 ( .B(n1094), .A(n1091), .S(n3136), .Y(n1105) );
  MUX2X1 U6846 ( .B(arr[1570]), .A(arr[1611]), .S(n2957), .Y(n1099) );
  MUX2X1 U6847 ( .B(arr[1488]), .A(arr[1529]), .S(n2957), .Y(n1098) );
  MUX2X1 U6848 ( .B(arr[1406]), .A(arr[1447]), .S(n2957), .Y(n1102) );
  MUX2X1 U6849 ( .B(arr[1324]), .A(arr[1365]), .S(n2957), .Y(n1101) );
  MUX2X1 U6850 ( .B(n1100), .A(n1097), .S(n3136), .Y(n1104) );
  MUX2X1 U6851 ( .B(n1103), .A(n1088), .S(n3182), .Y(n1137) );
  MUX2X1 U6852 ( .B(arr[1242]), .A(arr[1283]), .S(n2958), .Y(n1108) );
  MUX2X1 U6853 ( .B(arr[1160]), .A(arr[1201]), .S(n2958), .Y(n1107) );
  MUX2X1 U6854 ( .B(arr[1078]), .A(arr[1119]), .S(n2958), .Y(n1111) );
  MUX2X1 U6855 ( .B(arr[996]), .A(arr[1037]), .S(n2958), .Y(n1110) );
  MUX2X1 U6856 ( .B(n1109), .A(n1106), .S(n3137), .Y(n1120) );
  MUX2X1 U6857 ( .B(arr[914]), .A(arr[955]), .S(n2958), .Y(n1114) );
  MUX2X1 U6858 ( .B(arr[832]), .A(arr[873]), .S(n2958), .Y(n1113) );
  MUX2X1 U6859 ( .B(arr[750]), .A(arr[791]), .S(n2958), .Y(n1117) );
  MUX2X1 U6860 ( .B(arr[668]), .A(arr[709]), .S(n2958), .Y(n1116) );
  MUX2X1 U6861 ( .B(n1115), .A(n1112), .S(n3137), .Y(n1119) );
  MUX2X1 U6862 ( .B(arr[586]), .A(arr[627]), .S(n2958), .Y(n1123) );
  MUX2X1 U6863 ( .B(arr[504]), .A(arr[545]), .S(n2958), .Y(n1122) );
  MUX2X1 U6864 ( .B(arr[422]), .A(arr[463]), .S(n2958), .Y(n1126) );
  MUX2X1 U6865 ( .B(arr[340]), .A(arr[381]), .S(n2958), .Y(n1125) );
  MUX2X1 U6866 ( .B(n1124), .A(n1121), .S(n3137), .Y(n1135) );
  MUX2X1 U6867 ( .B(arr[258]), .A(arr[299]), .S(n2959), .Y(n1129) );
  MUX2X1 U6868 ( .B(arr[176]), .A(arr[217]), .S(n2959), .Y(n1128) );
  MUX2X1 U6869 ( .B(arr[94]), .A(arr[135]), .S(n2959), .Y(n1132) );
  MUX2X1 U6870 ( .B(arr[12]), .A(arr[53]), .S(n2959), .Y(n1131) );
  MUX2X1 U6871 ( .B(n1130), .A(n1127), .S(n3137), .Y(n1134) );
  MUX2X1 U6872 ( .B(n1133), .A(n1118), .S(n3182), .Y(n1136) );
  MUX2X1 U6873 ( .B(arr[2555]), .A(arr[2596]), .S(n2959), .Y(n1140) );
  MUX2X1 U6874 ( .B(arr[2473]), .A(arr[2514]), .S(n2959), .Y(n1139) );
  MUX2X1 U6875 ( .B(arr[2391]), .A(arr[2432]), .S(n2959), .Y(n1143) );
  MUX2X1 U6876 ( .B(arr[2309]), .A(arr[2350]), .S(n2959), .Y(n1142) );
  MUX2X1 U6877 ( .B(n1141), .A(n1138), .S(n3137), .Y(n1152) );
  MUX2X1 U6878 ( .B(arr[2227]), .A(arr[2268]), .S(n2959), .Y(n1146) );
  MUX2X1 U6879 ( .B(arr[2145]), .A(arr[2186]), .S(n2959), .Y(n1145) );
  MUX2X1 U6880 ( .B(arr[2063]), .A(arr[2104]), .S(n2959), .Y(n1149) );
  MUX2X1 U6881 ( .B(arr[1981]), .A(arr[2022]), .S(n2959), .Y(n1148) );
  MUX2X1 U6882 ( .B(n1147), .A(n1144), .S(n3137), .Y(n1151) );
  MUX2X1 U6883 ( .B(arr[1899]), .A(arr[1940]), .S(n2960), .Y(n1155) );
  MUX2X1 U6884 ( .B(arr[1817]), .A(arr[1858]), .S(n2960), .Y(n1154) );
  MUX2X1 U6885 ( .B(arr[1735]), .A(arr[1776]), .S(n2960), .Y(n1158) );
  MUX2X1 U6886 ( .B(arr[1653]), .A(arr[1694]), .S(n2960), .Y(n1157) );
  MUX2X1 U6887 ( .B(n1156), .A(n1153), .S(n3137), .Y(n1167) );
  MUX2X1 U6888 ( .B(arr[1571]), .A(arr[1612]), .S(n2960), .Y(n1161) );
  MUX2X1 U6889 ( .B(arr[1489]), .A(arr[1530]), .S(n2960), .Y(n1160) );
  MUX2X1 U6890 ( .B(arr[1407]), .A(arr[1448]), .S(n2960), .Y(n1164) );
  MUX2X1 U6891 ( .B(arr[1325]), .A(arr[1366]), .S(n2960), .Y(n1163) );
  MUX2X1 U6892 ( .B(n1162), .A(n1159), .S(n3137), .Y(n1166) );
  MUX2X1 U6893 ( .B(n1165), .A(n1150), .S(n3182), .Y(n1199) );
  MUX2X1 U6894 ( .B(arr[1243]), .A(arr[1284]), .S(n2960), .Y(n1170) );
  MUX2X1 U6895 ( .B(arr[1161]), .A(arr[1202]), .S(n2960), .Y(n1169) );
  MUX2X1 U6896 ( .B(arr[1079]), .A(arr[1120]), .S(n2960), .Y(n1173) );
  MUX2X1 U6897 ( .B(arr[997]), .A(arr[1038]), .S(n2960), .Y(n1172) );
  MUX2X1 U6898 ( .B(n1171), .A(n1168), .S(n3137), .Y(n1182) );
  MUX2X1 U6899 ( .B(arr[915]), .A(arr[956]), .S(n2961), .Y(n1176) );
  MUX2X1 U6900 ( .B(arr[833]), .A(arr[874]), .S(n2961), .Y(n1175) );
  MUX2X1 U6901 ( .B(arr[751]), .A(arr[792]), .S(n2961), .Y(n1179) );
  MUX2X1 U6902 ( .B(arr[669]), .A(arr[710]), .S(n2961), .Y(n1178) );
  MUX2X1 U6903 ( .B(n1177), .A(n1174), .S(n3137), .Y(n1181) );
  MUX2X1 U6904 ( .B(arr[587]), .A(arr[628]), .S(n2961), .Y(n1185) );
  MUX2X1 U6905 ( .B(arr[505]), .A(arr[546]), .S(n2961), .Y(n1184) );
  MUX2X1 U6906 ( .B(arr[423]), .A(arr[464]), .S(n2961), .Y(n1188) );
  MUX2X1 U6907 ( .B(arr[341]), .A(arr[382]), .S(n2961), .Y(n1187) );
  MUX2X1 U6908 ( .B(n1186), .A(n1183), .S(n3137), .Y(n1197) );
  MUX2X1 U6909 ( .B(arr[259]), .A(arr[300]), .S(n2961), .Y(n1191) );
  MUX2X1 U6910 ( .B(arr[177]), .A(arr[218]), .S(n2961), .Y(n1190) );
  MUX2X1 U6911 ( .B(arr[95]), .A(arr[136]), .S(n2961), .Y(n1194) );
  MUX2X1 U6912 ( .B(arr[13]), .A(arr[54]), .S(n2961), .Y(n1193) );
  MUX2X1 U6913 ( .B(n1192), .A(n1189), .S(n3137), .Y(n1196) );
  MUX2X1 U6914 ( .B(n1195), .A(n1180), .S(n3182), .Y(n1198) );
  MUX2X1 U6915 ( .B(arr[2556]), .A(arr[2597]), .S(n2962), .Y(n1202) );
  MUX2X1 U6916 ( .B(arr[2474]), .A(arr[2515]), .S(n2962), .Y(n1201) );
  MUX2X1 U6917 ( .B(arr[2392]), .A(arr[2433]), .S(n2962), .Y(n1205) );
  MUX2X1 U6918 ( .B(arr[2310]), .A(arr[2351]), .S(n2962), .Y(n1204) );
  MUX2X1 U6919 ( .B(n1203), .A(n1200), .S(n3138), .Y(n1214) );
  MUX2X1 U6920 ( .B(arr[2228]), .A(arr[2269]), .S(n2962), .Y(n1208) );
  MUX2X1 U6921 ( .B(arr[2146]), .A(arr[2187]), .S(n2962), .Y(n1207) );
  MUX2X1 U6922 ( .B(arr[2064]), .A(arr[2105]), .S(n2962), .Y(n1211) );
  MUX2X1 U6923 ( .B(arr[1982]), .A(arr[2023]), .S(n2962), .Y(n1210) );
  MUX2X1 U6924 ( .B(n1209), .A(n1206), .S(n3138), .Y(n1213) );
  MUX2X1 U6925 ( .B(arr[1900]), .A(arr[1941]), .S(n2962), .Y(n1217) );
  MUX2X1 U6926 ( .B(arr[1818]), .A(arr[1859]), .S(n2962), .Y(n1216) );
  MUX2X1 U6927 ( .B(arr[1736]), .A(arr[1777]), .S(n2962), .Y(n1220) );
  MUX2X1 U6928 ( .B(arr[1654]), .A(arr[1695]), .S(n2962), .Y(n1219) );
  MUX2X1 U6929 ( .B(n1218), .A(n1215), .S(n3138), .Y(n1229) );
  MUX2X1 U6930 ( .B(arr[1572]), .A(arr[1613]), .S(n2963), .Y(n1223) );
  MUX2X1 U6931 ( .B(arr[1490]), .A(arr[1531]), .S(n2963), .Y(n1222) );
  MUX2X1 U6932 ( .B(arr[1408]), .A(arr[1449]), .S(n2963), .Y(n1226) );
  MUX2X1 U6933 ( .B(arr[1326]), .A(arr[1367]), .S(n2963), .Y(n1225) );
  MUX2X1 U6934 ( .B(n1224), .A(n1221), .S(n3138), .Y(n1228) );
  MUX2X1 U6935 ( .B(n1227), .A(n1212), .S(n3182), .Y(n1261) );
  MUX2X1 U6936 ( .B(arr[1244]), .A(arr[1285]), .S(n2963), .Y(n1232) );
  MUX2X1 U6937 ( .B(arr[1162]), .A(arr[1203]), .S(n2963), .Y(n1231) );
  MUX2X1 U6938 ( .B(arr[1080]), .A(arr[1121]), .S(n2963), .Y(n1235) );
  MUX2X1 U6939 ( .B(arr[998]), .A(arr[1039]), .S(n2963), .Y(n1234) );
  MUX2X1 U6940 ( .B(n1233), .A(n1230), .S(n3138), .Y(n1244) );
  MUX2X1 U6941 ( .B(arr[916]), .A(arr[957]), .S(n2963), .Y(n1238) );
  MUX2X1 U6942 ( .B(arr[834]), .A(arr[875]), .S(n2963), .Y(n1237) );
  MUX2X1 U6943 ( .B(arr[752]), .A(arr[793]), .S(n2963), .Y(n1241) );
  MUX2X1 U6944 ( .B(arr[670]), .A(arr[711]), .S(n2963), .Y(n1240) );
  MUX2X1 U6945 ( .B(n1239), .A(n1236), .S(n3138), .Y(n1243) );
  MUX2X1 U6946 ( .B(arr[588]), .A(arr[629]), .S(n2964), .Y(n1247) );
  MUX2X1 U6947 ( .B(arr[506]), .A(arr[547]), .S(n2964), .Y(n1246) );
  MUX2X1 U6948 ( .B(arr[424]), .A(arr[465]), .S(n2964), .Y(n1250) );
  MUX2X1 U6949 ( .B(arr[342]), .A(arr[383]), .S(n2964), .Y(n1249) );
  MUX2X1 U6950 ( .B(n1248), .A(n1245), .S(n3138), .Y(n1259) );
  MUX2X1 U6951 ( .B(arr[260]), .A(arr[301]), .S(n2964), .Y(n1253) );
  MUX2X1 U6952 ( .B(arr[178]), .A(arr[219]), .S(n2964), .Y(n1252) );
  MUX2X1 U6953 ( .B(arr[96]), .A(arr[137]), .S(n2964), .Y(n1256) );
  MUX2X1 U6954 ( .B(arr[14]), .A(arr[55]), .S(n2964), .Y(n1255) );
  MUX2X1 U6955 ( .B(n1254), .A(n1251), .S(n3138), .Y(n1258) );
  MUX2X1 U6956 ( .B(n1257), .A(n1242), .S(n3182), .Y(n1260) );
  MUX2X1 U6957 ( .B(arr[2557]), .A(arr[2598]), .S(n2964), .Y(n1264) );
  MUX2X1 U6958 ( .B(arr[2475]), .A(arr[2516]), .S(n2964), .Y(n1263) );
  MUX2X1 U6959 ( .B(arr[2393]), .A(arr[2434]), .S(n2964), .Y(n1267) );
  MUX2X1 U6960 ( .B(arr[2311]), .A(arr[2352]), .S(n2964), .Y(n1266) );
  MUX2X1 U6961 ( .B(n1265), .A(n1262), .S(n3138), .Y(n1276) );
  MUX2X1 U6962 ( .B(arr[2229]), .A(arr[2270]), .S(n2965), .Y(n1270) );
  MUX2X1 U6963 ( .B(arr[2147]), .A(arr[2188]), .S(n2965), .Y(n1269) );
  MUX2X1 U6964 ( .B(arr[2065]), .A(arr[2106]), .S(n2965), .Y(n1273) );
  MUX2X1 U6965 ( .B(arr[1983]), .A(arr[2024]), .S(n2965), .Y(n1272) );
  MUX2X1 U6966 ( .B(n1271), .A(n1268), .S(n3138), .Y(n1275) );
  MUX2X1 U6967 ( .B(arr[1901]), .A(arr[1942]), .S(n2965), .Y(n1279) );
  MUX2X1 U6968 ( .B(arr[1819]), .A(arr[1860]), .S(n2965), .Y(n1278) );
  MUX2X1 U6969 ( .B(arr[1737]), .A(arr[1778]), .S(n2965), .Y(n1282) );
  MUX2X1 U6970 ( .B(arr[1655]), .A(arr[1696]), .S(n2965), .Y(n1281) );
  MUX2X1 U6971 ( .B(n1280), .A(n1277), .S(n3138), .Y(n1291) );
  MUX2X1 U6972 ( .B(arr[1573]), .A(arr[1614]), .S(n2965), .Y(n1285) );
  MUX2X1 U6973 ( .B(arr[1491]), .A(arr[1532]), .S(n2965), .Y(n1284) );
  MUX2X1 U6974 ( .B(arr[1409]), .A(arr[1450]), .S(n2965), .Y(n1288) );
  MUX2X1 U6975 ( .B(arr[1327]), .A(arr[1368]), .S(n2965), .Y(n1287) );
  MUX2X1 U6976 ( .B(n1286), .A(n1283), .S(n3138), .Y(n1290) );
  MUX2X1 U6977 ( .B(n1289), .A(n1274), .S(n3182), .Y(n1323) );
  MUX2X1 U6978 ( .B(arr[1245]), .A(arr[1286]), .S(n2966), .Y(n1294) );
  MUX2X1 U6979 ( .B(arr[1163]), .A(arr[1204]), .S(n2966), .Y(n1293) );
  MUX2X1 U6980 ( .B(arr[1081]), .A(arr[1122]), .S(n2966), .Y(n1297) );
  MUX2X1 U6981 ( .B(arr[999]), .A(arr[1040]), .S(n2966), .Y(n1296) );
  MUX2X1 U6982 ( .B(n1295), .A(n1292), .S(n3139), .Y(n1306) );
  MUX2X1 U6983 ( .B(arr[917]), .A(arr[958]), .S(n2966), .Y(n1300) );
  MUX2X1 U6984 ( .B(arr[835]), .A(arr[876]), .S(n2966), .Y(n1299) );
  MUX2X1 U6985 ( .B(arr[753]), .A(arr[794]), .S(n2966), .Y(n1303) );
  MUX2X1 U6986 ( .B(arr[671]), .A(arr[712]), .S(n2966), .Y(n1302) );
  MUX2X1 U6987 ( .B(n1301), .A(n1298), .S(n3139), .Y(n1305) );
  MUX2X1 U6988 ( .B(arr[589]), .A(arr[630]), .S(n2966), .Y(n1309) );
  MUX2X1 U6989 ( .B(arr[507]), .A(arr[548]), .S(n2966), .Y(n1308) );
  MUX2X1 U6990 ( .B(arr[425]), .A(arr[466]), .S(n2966), .Y(n1312) );
  MUX2X1 U6991 ( .B(arr[343]), .A(arr[384]), .S(n2966), .Y(n1311) );
  MUX2X1 U6992 ( .B(n1310), .A(n1307), .S(n3139), .Y(n1321) );
  MUX2X1 U6993 ( .B(arr[261]), .A(arr[302]), .S(n2967), .Y(n1315) );
  MUX2X1 U6994 ( .B(arr[179]), .A(arr[220]), .S(n2967), .Y(n1314) );
  MUX2X1 U6995 ( .B(arr[97]), .A(arr[138]), .S(n2967), .Y(n1318) );
  MUX2X1 U6996 ( .B(arr[15]), .A(arr[56]), .S(n2967), .Y(n1317) );
  MUX2X1 U6997 ( .B(n1316), .A(n1313), .S(n3139), .Y(n1320) );
  MUX2X1 U6998 ( .B(n1319), .A(n1304), .S(n3182), .Y(n1322) );
  MUX2X1 U6999 ( .B(arr[2558]), .A(arr[2599]), .S(n2967), .Y(n1326) );
  MUX2X1 U7000 ( .B(arr[2476]), .A(arr[2517]), .S(n2967), .Y(n1325) );
  MUX2X1 U7001 ( .B(arr[2394]), .A(arr[2435]), .S(n2967), .Y(n1329) );
  MUX2X1 U7002 ( .B(arr[2312]), .A(arr[2353]), .S(n2967), .Y(n1328) );
  MUX2X1 U7003 ( .B(n1327), .A(n1324), .S(n3139), .Y(n1338) );
  MUX2X1 U7004 ( .B(arr[2230]), .A(arr[2271]), .S(n2967), .Y(n1332) );
  MUX2X1 U7005 ( .B(arr[2148]), .A(arr[2189]), .S(n2967), .Y(n1331) );
  MUX2X1 U7006 ( .B(arr[2066]), .A(arr[2107]), .S(n2967), .Y(n1335) );
  MUX2X1 U7007 ( .B(arr[1984]), .A(arr[2025]), .S(n2967), .Y(n1334) );
  MUX2X1 U7008 ( .B(n1333), .A(n1330), .S(n3139), .Y(n1337) );
  MUX2X1 U7009 ( .B(arr[1902]), .A(arr[1943]), .S(n2968), .Y(n1341) );
  MUX2X1 U7010 ( .B(arr[1820]), .A(arr[1861]), .S(n2968), .Y(n1340) );
  MUX2X1 U7011 ( .B(arr[1738]), .A(arr[1779]), .S(n2968), .Y(n1344) );
  MUX2X1 U7012 ( .B(arr[1656]), .A(arr[1697]), .S(n2968), .Y(n1343) );
  MUX2X1 U7013 ( .B(n1342), .A(n1339), .S(n3139), .Y(n1353) );
  MUX2X1 U7014 ( .B(arr[1574]), .A(arr[1615]), .S(n2968), .Y(n1347) );
  MUX2X1 U7015 ( .B(arr[1492]), .A(arr[1533]), .S(n2968), .Y(n1346) );
  MUX2X1 U7016 ( .B(arr[1410]), .A(arr[1451]), .S(n2968), .Y(n1350) );
  MUX2X1 U7017 ( .B(arr[1328]), .A(arr[1369]), .S(n2968), .Y(n1349) );
  MUX2X1 U7018 ( .B(n1348), .A(n1345), .S(n3139), .Y(n1352) );
  MUX2X1 U7019 ( .B(n1351), .A(n1336), .S(n3182), .Y(n1385) );
  MUX2X1 U7020 ( .B(arr[1246]), .A(arr[1287]), .S(n2968), .Y(n1356) );
  MUX2X1 U7021 ( .B(arr[1164]), .A(arr[1205]), .S(n2968), .Y(n1355) );
  MUX2X1 U7022 ( .B(arr[1082]), .A(arr[1123]), .S(n2968), .Y(n1359) );
  MUX2X1 U7023 ( .B(arr[1000]), .A(arr[1041]), .S(n2968), .Y(n1358) );
  MUX2X1 U7024 ( .B(n1357), .A(n1354), .S(n3139), .Y(n1368) );
  MUX2X1 U7025 ( .B(arr[918]), .A(arr[959]), .S(n2969), .Y(n1362) );
  MUX2X1 U7026 ( .B(arr[836]), .A(arr[877]), .S(n2969), .Y(n1361) );
  MUX2X1 U7027 ( .B(arr[754]), .A(arr[795]), .S(n2969), .Y(n1365) );
  MUX2X1 U7028 ( .B(arr[672]), .A(arr[713]), .S(n2969), .Y(n1364) );
  MUX2X1 U7029 ( .B(n1363), .A(n1360), .S(n3139), .Y(n1367) );
  MUX2X1 U7030 ( .B(arr[590]), .A(arr[631]), .S(n2969), .Y(n1371) );
  MUX2X1 U7031 ( .B(arr[508]), .A(arr[549]), .S(n2969), .Y(n1370) );
  MUX2X1 U7032 ( .B(arr[426]), .A(arr[467]), .S(n2969), .Y(n1374) );
  MUX2X1 U7033 ( .B(arr[344]), .A(arr[385]), .S(n2969), .Y(n1373) );
  MUX2X1 U7034 ( .B(n1372), .A(n1369), .S(n3139), .Y(n1383) );
  MUX2X1 U7035 ( .B(arr[262]), .A(arr[303]), .S(n2969), .Y(n1377) );
  MUX2X1 U7036 ( .B(arr[180]), .A(arr[221]), .S(n2969), .Y(n1376) );
  MUX2X1 U7037 ( .B(arr[98]), .A(arr[139]), .S(n2969), .Y(n1380) );
  MUX2X1 U7038 ( .B(arr[16]), .A(arr[57]), .S(n2969), .Y(n1379) );
  MUX2X1 U7039 ( .B(n1378), .A(n1375), .S(n3139), .Y(n1382) );
  MUX2X1 U7040 ( .B(n1381), .A(n1366), .S(n3182), .Y(n1384) );
  MUX2X1 U7041 ( .B(arr[2559]), .A(arr[2600]), .S(n2970), .Y(n1388) );
  MUX2X1 U7042 ( .B(arr[2477]), .A(arr[2518]), .S(n2970), .Y(n1387) );
  MUX2X1 U7043 ( .B(arr[2395]), .A(arr[2436]), .S(n2970), .Y(n1391) );
  MUX2X1 U7044 ( .B(arr[2313]), .A(arr[2354]), .S(n2970), .Y(n1390) );
  MUX2X1 U7045 ( .B(n1389), .A(n1386), .S(n3140), .Y(n1400) );
  MUX2X1 U7046 ( .B(arr[2231]), .A(arr[2272]), .S(n2970), .Y(n1394) );
  MUX2X1 U7047 ( .B(arr[2149]), .A(arr[2190]), .S(n2970), .Y(n1393) );
  MUX2X1 U7048 ( .B(arr[2067]), .A(arr[2108]), .S(n2970), .Y(n1397) );
  MUX2X1 U7049 ( .B(arr[1985]), .A(arr[2026]), .S(n2970), .Y(n1396) );
  MUX2X1 U7050 ( .B(n1395), .A(n1392), .S(n3140), .Y(n1399) );
  MUX2X1 U7051 ( .B(arr[1903]), .A(arr[1944]), .S(n2970), .Y(n1403) );
  MUX2X1 U7052 ( .B(arr[1821]), .A(arr[1862]), .S(n2970), .Y(n1402) );
  MUX2X1 U7053 ( .B(arr[1739]), .A(arr[1780]), .S(n2970), .Y(n1406) );
  MUX2X1 U7054 ( .B(arr[1657]), .A(arr[1698]), .S(n2970), .Y(n1405) );
  MUX2X1 U7055 ( .B(n1404), .A(n1401), .S(n3140), .Y(n1415) );
  MUX2X1 U7056 ( .B(arr[1575]), .A(arr[1616]), .S(n2971), .Y(n1409) );
  MUX2X1 U7057 ( .B(arr[1493]), .A(arr[1534]), .S(n2971), .Y(n1408) );
  MUX2X1 U7058 ( .B(arr[1411]), .A(arr[1452]), .S(n2971), .Y(n1412) );
  MUX2X1 U7059 ( .B(arr[1329]), .A(arr[1370]), .S(n2971), .Y(n1411) );
  MUX2X1 U7060 ( .B(n1410), .A(n1407), .S(n3140), .Y(n1414) );
  MUX2X1 U7061 ( .B(n1413), .A(n1398), .S(n3183), .Y(n1447) );
  MUX2X1 U7062 ( .B(arr[1247]), .A(arr[1288]), .S(n2971), .Y(n1418) );
  MUX2X1 U7063 ( .B(arr[1165]), .A(arr[1206]), .S(n2971), .Y(n1417) );
  MUX2X1 U7064 ( .B(arr[1083]), .A(arr[1124]), .S(n2971), .Y(n1421) );
  MUX2X1 U7065 ( .B(arr[1001]), .A(arr[1042]), .S(n2971), .Y(n1420) );
  MUX2X1 U7066 ( .B(n1419), .A(n1416), .S(n3140), .Y(n1430) );
  MUX2X1 U7067 ( .B(arr[919]), .A(arr[960]), .S(n2971), .Y(n1424) );
  MUX2X1 U7068 ( .B(arr[837]), .A(arr[878]), .S(n2971), .Y(n1423) );
  MUX2X1 U7069 ( .B(arr[755]), .A(arr[796]), .S(n2971), .Y(n1427) );
  MUX2X1 U7070 ( .B(arr[673]), .A(arr[714]), .S(n2971), .Y(n1426) );
  MUX2X1 U7071 ( .B(n1425), .A(n1422), .S(n3140), .Y(n1429) );
  MUX2X1 U7072 ( .B(arr[591]), .A(arr[632]), .S(n2972), .Y(n1433) );
  MUX2X1 U7073 ( .B(arr[509]), .A(arr[550]), .S(n2972), .Y(n1432) );
  MUX2X1 U7074 ( .B(arr[427]), .A(arr[468]), .S(n2972), .Y(n1436) );
  MUX2X1 U7075 ( .B(arr[345]), .A(arr[386]), .S(n2972), .Y(n1435) );
  MUX2X1 U7076 ( .B(n1434), .A(n1431), .S(n3140), .Y(n1445) );
  MUX2X1 U7077 ( .B(arr[263]), .A(arr[304]), .S(n2972), .Y(n1439) );
  MUX2X1 U7078 ( .B(arr[181]), .A(arr[222]), .S(n2972), .Y(n1438) );
  MUX2X1 U7079 ( .B(arr[99]), .A(arr[140]), .S(n2972), .Y(n1442) );
  MUX2X1 U7080 ( .B(arr[17]), .A(arr[58]), .S(n2972), .Y(n1441) );
  MUX2X1 U7081 ( .B(n1440), .A(n1437), .S(n3140), .Y(n1444) );
  MUX2X1 U7082 ( .B(n1443), .A(n1428), .S(n3183), .Y(n1446) );
  MUX2X1 U7083 ( .B(arr[2560]), .A(arr[2601]), .S(n2972), .Y(n1450) );
  MUX2X1 U7084 ( .B(arr[2478]), .A(arr[2519]), .S(n2972), .Y(n1449) );
  MUX2X1 U7085 ( .B(arr[2396]), .A(arr[2437]), .S(n2972), .Y(n1453) );
  MUX2X1 U7086 ( .B(arr[2314]), .A(arr[2355]), .S(n2972), .Y(n1452) );
  MUX2X1 U7087 ( .B(n1451), .A(n1448), .S(n3140), .Y(n1462) );
  MUX2X1 U7088 ( .B(arr[2232]), .A(arr[2273]), .S(n2973), .Y(n1456) );
  MUX2X1 U7089 ( .B(arr[2150]), .A(arr[2191]), .S(n2973), .Y(n1455) );
  MUX2X1 U7090 ( .B(arr[2068]), .A(arr[2109]), .S(n2973), .Y(n1459) );
  MUX2X1 U7091 ( .B(arr[1986]), .A(arr[2027]), .S(n2973), .Y(n1458) );
  MUX2X1 U7092 ( .B(n1457), .A(n1454), .S(n3140), .Y(n1461) );
  MUX2X1 U7093 ( .B(arr[1904]), .A(arr[1945]), .S(n2973), .Y(n1465) );
  MUX2X1 U7094 ( .B(arr[1822]), .A(arr[1863]), .S(n2973), .Y(n1464) );
  MUX2X1 U7095 ( .B(arr[1740]), .A(arr[1781]), .S(n2973), .Y(n1468) );
  MUX2X1 U7096 ( .B(arr[1658]), .A(arr[1699]), .S(n2973), .Y(n1467) );
  MUX2X1 U7097 ( .B(n1466), .A(n1463), .S(n3140), .Y(n1477) );
  MUX2X1 U7098 ( .B(arr[1576]), .A(arr[1617]), .S(n2973), .Y(n1471) );
  MUX2X1 U7099 ( .B(arr[1494]), .A(arr[1535]), .S(n2973), .Y(n1470) );
  MUX2X1 U7100 ( .B(arr[1412]), .A(arr[1453]), .S(n2973), .Y(n1474) );
  MUX2X1 U7101 ( .B(arr[1330]), .A(arr[1371]), .S(n2973), .Y(n1473) );
  MUX2X1 U7102 ( .B(n1472), .A(n1469), .S(n3140), .Y(n1476) );
  MUX2X1 U7103 ( .B(n1475), .A(n1460), .S(n3183), .Y(n1509) );
  MUX2X1 U7104 ( .B(arr[1248]), .A(arr[1289]), .S(n2974), .Y(n1480) );
  MUX2X1 U7105 ( .B(arr[1166]), .A(arr[1207]), .S(n2974), .Y(n1479) );
  MUX2X1 U7106 ( .B(arr[1084]), .A(arr[1125]), .S(n2974), .Y(n1483) );
  MUX2X1 U7107 ( .B(arr[1002]), .A(arr[1043]), .S(n2974), .Y(n1482) );
  MUX2X1 U7108 ( .B(n1481), .A(n1478), .S(n3141), .Y(n1492) );
  MUX2X1 U7109 ( .B(arr[920]), .A(arr[961]), .S(n2974), .Y(n1486) );
  MUX2X1 U7110 ( .B(arr[838]), .A(arr[879]), .S(n2974), .Y(n1485) );
  MUX2X1 U7111 ( .B(arr[756]), .A(arr[797]), .S(n2974), .Y(n1489) );
  MUX2X1 U7112 ( .B(arr[674]), .A(arr[715]), .S(n2974), .Y(n1488) );
  MUX2X1 U7113 ( .B(n1487), .A(n1484), .S(n3141), .Y(n1491) );
  MUX2X1 U7114 ( .B(arr[592]), .A(arr[633]), .S(n2974), .Y(n1495) );
  MUX2X1 U7115 ( .B(arr[510]), .A(arr[551]), .S(n2974), .Y(n1494) );
  MUX2X1 U7116 ( .B(arr[428]), .A(arr[469]), .S(n2974), .Y(n1498) );
  MUX2X1 U7117 ( .B(arr[346]), .A(arr[387]), .S(n2974), .Y(n1497) );
  MUX2X1 U7118 ( .B(n1496), .A(n1493), .S(n3141), .Y(n1507) );
  MUX2X1 U7119 ( .B(arr[264]), .A(arr[305]), .S(n2975), .Y(n1501) );
  MUX2X1 U7120 ( .B(arr[182]), .A(arr[223]), .S(n2975), .Y(n1500) );
  MUX2X1 U7121 ( .B(arr[100]), .A(arr[141]), .S(n2975), .Y(n1504) );
  MUX2X1 U7122 ( .B(arr[18]), .A(arr[59]), .S(n2975), .Y(n1503) );
  MUX2X1 U7123 ( .B(n1502), .A(n1499), .S(n3141), .Y(n1506) );
  MUX2X1 U7124 ( .B(n1505), .A(n1490), .S(n3183), .Y(n1508) );
  MUX2X1 U7125 ( .B(arr[2561]), .A(arr[2602]), .S(n2975), .Y(n1512) );
  MUX2X1 U7126 ( .B(arr[2479]), .A(arr[2520]), .S(n2975), .Y(n1511) );
  MUX2X1 U7127 ( .B(arr[2397]), .A(arr[2438]), .S(n2975), .Y(n1515) );
  MUX2X1 U7128 ( .B(arr[2315]), .A(arr[2356]), .S(n2975), .Y(n1514) );
  MUX2X1 U7129 ( .B(n1513), .A(n1510), .S(n3141), .Y(n1524) );
  MUX2X1 U7130 ( .B(arr[2233]), .A(arr[2274]), .S(n2975), .Y(n1518) );
  MUX2X1 U7131 ( .B(arr[2151]), .A(arr[2192]), .S(n2975), .Y(n1517) );
  MUX2X1 U7132 ( .B(arr[2069]), .A(arr[2110]), .S(n2975), .Y(n1521) );
  MUX2X1 U7133 ( .B(arr[1987]), .A(arr[2028]), .S(n2975), .Y(n1520) );
  MUX2X1 U7134 ( .B(n1519), .A(n1516), .S(n3141), .Y(n1523) );
  MUX2X1 U7135 ( .B(arr[1905]), .A(arr[1946]), .S(n2976), .Y(n1527) );
  MUX2X1 U7136 ( .B(arr[1823]), .A(arr[1864]), .S(n2976), .Y(n1526) );
  MUX2X1 U7137 ( .B(arr[1741]), .A(arr[1782]), .S(n2976), .Y(n1530) );
  MUX2X1 U7138 ( .B(arr[1659]), .A(arr[1700]), .S(n2976), .Y(n1529) );
  MUX2X1 U7139 ( .B(n1528), .A(n1525), .S(n3141), .Y(n1539) );
  MUX2X1 U7140 ( .B(arr[1577]), .A(arr[1618]), .S(n2976), .Y(n1533) );
  MUX2X1 U7141 ( .B(arr[1495]), .A(arr[1536]), .S(n2976), .Y(n1532) );
  MUX2X1 U7142 ( .B(arr[1413]), .A(arr[1454]), .S(n2976), .Y(n1536) );
  MUX2X1 U7143 ( .B(arr[1331]), .A(arr[1372]), .S(n2976), .Y(n1535) );
  MUX2X1 U7144 ( .B(n1534), .A(n1531), .S(n3141), .Y(n1538) );
  MUX2X1 U7145 ( .B(n1537), .A(n1522), .S(n3183), .Y(n1571) );
  MUX2X1 U7146 ( .B(arr[1249]), .A(arr[1290]), .S(n2976), .Y(n1542) );
  MUX2X1 U7147 ( .B(arr[1167]), .A(arr[1208]), .S(n2976), .Y(n1541) );
  MUX2X1 U7148 ( .B(arr[1085]), .A(arr[1126]), .S(n2976), .Y(n1545) );
  MUX2X1 U7149 ( .B(arr[1003]), .A(arr[1044]), .S(n2976), .Y(n1544) );
  MUX2X1 U7150 ( .B(n1543), .A(n1540), .S(n3141), .Y(n1554) );
  MUX2X1 U7151 ( .B(arr[921]), .A(arr[962]), .S(n2977), .Y(n1548) );
  MUX2X1 U7152 ( .B(arr[839]), .A(arr[880]), .S(n2977), .Y(n1547) );
  MUX2X1 U7153 ( .B(arr[757]), .A(arr[798]), .S(n2977), .Y(n1551) );
  MUX2X1 U7154 ( .B(arr[675]), .A(arr[716]), .S(n2977), .Y(n1550) );
  MUX2X1 U7155 ( .B(n1549), .A(n1546), .S(n3141), .Y(n1553) );
  MUX2X1 U7156 ( .B(arr[593]), .A(arr[634]), .S(n2977), .Y(n1557) );
  MUX2X1 U7157 ( .B(arr[511]), .A(arr[552]), .S(n2977), .Y(n1556) );
  MUX2X1 U7158 ( .B(arr[429]), .A(arr[470]), .S(n2977), .Y(n1560) );
  MUX2X1 U7159 ( .B(arr[347]), .A(arr[388]), .S(n2977), .Y(n1559) );
  MUX2X1 U7160 ( .B(n1558), .A(n1555), .S(n3141), .Y(n1569) );
  MUX2X1 U7161 ( .B(arr[265]), .A(arr[306]), .S(n2977), .Y(n1563) );
  MUX2X1 U7162 ( .B(arr[183]), .A(arr[224]), .S(n2977), .Y(n1562) );
  MUX2X1 U7163 ( .B(arr[101]), .A(arr[142]), .S(n2977), .Y(n1566) );
  MUX2X1 U7164 ( .B(arr[19]), .A(arr[60]), .S(n2977), .Y(n1565) );
  MUX2X1 U7165 ( .B(n1564), .A(n1561), .S(n3141), .Y(n1568) );
  MUX2X1 U7166 ( .B(n1567), .A(n1552), .S(n3183), .Y(n1570) );
  MUX2X1 U7167 ( .B(arr[2562]), .A(arr[2603]), .S(n2978), .Y(n1574) );
  MUX2X1 U7168 ( .B(arr[2480]), .A(arr[2521]), .S(n2978), .Y(n1573) );
  MUX2X1 U7169 ( .B(arr[2398]), .A(arr[2439]), .S(n2978), .Y(n1577) );
  MUX2X1 U7170 ( .B(arr[2316]), .A(arr[2357]), .S(n2978), .Y(n1576) );
  MUX2X1 U7171 ( .B(n1575), .A(n1572), .S(n3142), .Y(n1586) );
  MUX2X1 U7172 ( .B(arr[2234]), .A(arr[2275]), .S(n2978), .Y(n1580) );
  MUX2X1 U7173 ( .B(arr[2152]), .A(arr[2193]), .S(n2978), .Y(n1579) );
  MUX2X1 U7174 ( .B(arr[2070]), .A(arr[2111]), .S(n2978), .Y(n1583) );
  MUX2X1 U7175 ( .B(arr[1988]), .A(arr[2029]), .S(n2978), .Y(n1582) );
  MUX2X1 U7176 ( .B(n1581), .A(n1578), .S(n3142), .Y(n1585) );
  MUX2X1 U7177 ( .B(arr[1906]), .A(arr[1947]), .S(n2978), .Y(n1589) );
  MUX2X1 U7178 ( .B(arr[1824]), .A(arr[1865]), .S(n2978), .Y(n1588) );
  MUX2X1 U7179 ( .B(arr[1742]), .A(arr[1783]), .S(n2978), .Y(n1592) );
  MUX2X1 U7180 ( .B(arr[1660]), .A(arr[1701]), .S(n2978), .Y(n1591) );
  MUX2X1 U7181 ( .B(n1590), .A(n1587), .S(n3142), .Y(n1601) );
  MUX2X1 U7182 ( .B(arr[1578]), .A(arr[1619]), .S(n2979), .Y(n1595) );
  MUX2X1 U7183 ( .B(arr[1496]), .A(arr[1537]), .S(n2979), .Y(n1594) );
  MUX2X1 U7184 ( .B(arr[1414]), .A(arr[1455]), .S(n2979), .Y(n1598) );
  MUX2X1 U7185 ( .B(arr[1332]), .A(arr[1373]), .S(n2979), .Y(n1597) );
  MUX2X1 U7186 ( .B(n1596), .A(n1593), .S(n3142), .Y(n1600) );
  MUX2X1 U7187 ( .B(n1599), .A(n1584), .S(n3183), .Y(n1633) );
  MUX2X1 U7188 ( .B(arr[1250]), .A(arr[1291]), .S(n2979), .Y(n1604) );
  MUX2X1 U7189 ( .B(arr[1168]), .A(arr[1209]), .S(n2979), .Y(n1603) );
  MUX2X1 U7190 ( .B(arr[1086]), .A(arr[1127]), .S(n2979), .Y(n1607) );
  MUX2X1 U7191 ( .B(arr[1004]), .A(arr[1045]), .S(n2979), .Y(n1606) );
  MUX2X1 U7192 ( .B(n1605), .A(n1602), .S(n3142), .Y(n1616) );
  MUX2X1 U7193 ( .B(arr[922]), .A(arr[963]), .S(n2979), .Y(n1610) );
  MUX2X1 U7194 ( .B(arr[840]), .A(arr[881]), .S(n2979), .Y(n1609) );
  MUX2X1 U7195 ( .B(arr[758]), .A(arr[799]), .S(n2979), .Y(n1613) );
  MUX2X1 U7196 ( .B(arr[676]), .A(arr[717]), .S(n2979), .Y(n1612) );
  MUX2X1 U7197 ( .B(n1611), .A(n1608), .S(n3142), .Y(n1615) );
  MUX2X1 U7198 ( .B(arr[594]), .A(arr[635]), .S(n2980), .Y(n1619) );
  MUX2X1 U7199 ( .B(arr[512]), .A(arr[553]), .S(n2980), .Y(n1618) );
  MUX2X1 U7200 ( .B(arr[430]), .A(arr[471]), .S(n2980), .Y(n1622) );
  MUX2X1 U7201 ( .B(arr[348]), .A(arr[389]), .S(n2980), .Y(n1621) );
  MUX2X1 U7202 ( .B(n1620), .A(n1617), .S(n3142), .Y(n1631) );
  MUX2X1 U7203 ( .B(arr[266]), .A(arr[307]), .S(n2980), .Y(n1625) );
  MUX2X1 U7204 ( .B(arr[184]), .A(arr[225]), .S(n2980), .Y(n1624) );
  MUX2X1 U7205 ( .B(arr[102]), .A(arr[143]), .S(n2980), .Y(n1628) );
  MUX2X1 U7206 ( .B(arr[20]), .A(arr[61]), .S(n2980), .Y(n1627) );
  MUX2X1 U7207 ( .B(n1626), .A(n1623), .S(n3142), .Y(n1630) );
  MUX2X1 U7208 ( .B(n1629), .A(n1614), .S(n3183), .Y(n1632) );
  MUX2X1 U7209 ( .B(arr[2563]), .A(arr[2604]), .S(n2980), .Y(n1636) );
  MUX2X1 U7210 ( .B(arr[2481]), .A(arr[2522]), .S(n2980), .Y(n1635) );
  MUX2X1 U7211 ( .B(arr[2399]), .A(arr[2440]), .S(n2980), .Y(n1639) );
  MUX2X1 U7212 ( .B(arr[2317]), .A(arr[2358]), .S(n2980), .Y(n1638) );
  MUX2X1 U7213 ( .B(n1637), .A(n1634), .S(n3142), .Y(n1648) );
  MUX2X1 U7214 ( .B(arr[2235]), .A(arr[2276]), .S(n2981), .Y(n1642) );
  MUX2X1 U7215 ( .B(arr[2153]), .A(arr[2194]), .S(n2981), .Y(n1641) );
  MUX2X1 U7216 ( .B(arr[2071]), .A(arr[2112]), .S(n2981), .Y(n1645) );
  MUX2X1 U7217 ( .B(arr[1989]), .A(arr[2030]), .S(n2981), .Y(n1644) );
  MUX2X1 U7218 ( .B(n1643), .A(n1640), .S(n3142), .Y(n1647) );
  MUX2X1 U7219 ( .B(arr[1907]), .A(arr[1948]), .S(n2981), .Y(n1651) );
  MUX2X1 U7220 ( .B(arr[1825]), .A(arr[1866]), .S(n2981), .Y(n1650) );
  MUX2X1 U7221 ( .B(arr[1743]), .A(arr[1784]), .S(n2981), .Y(n1654) );
  MUX2X1 U7222 ( .B(arr[1661]), .A(arr[1702]), .S(n2981), .Y(n1653) );
  MUX2X1 U7223 ( .B(n1652), .A(n1649), .S(n3142), .Y(n1663) );
  MUX2X1 U7224 ( .B(arr[1579]), .A(arr[1620]), .S(n2981), .Y(n1657) );
  MUX2X1 U7225 ( .B(arr[1497]), .A(arr[1538]), .S(n2981), .Y(n1656) );
  MUX2X1 U7226 ( .B(arr[1415]), .A(arr[1456]), .S(n2981), .Y(n1660) );
  MUX2X1 U7227 ( .B(arr[1333]), .A(arr[1374]), .S(n2981), .Y(n1659) );
  MUX2X1 U7228 ( .B(n1658), .A(n1655), .S(n3142), .Y(n1662) );
  MUX2X1 U7229 ( .B(n1661), .A(n1646), .S(n3183), .Y(n1695) );
  MUX2X1 U7230 ( .B(arr[1251]), .A(arr[1292]), .S(n2982), .Y(n1666) );
  MUX2X1 U7231 ( .B(arr[1169]), .A(arr[1210]), .S(n2982), .Y(n1665) );
  MUX2X1 U7232 ( .B(arr[1087]), .A(arr[1128]), .S(n2982), .Y(n1669) );
  MUX2X1 U7233 ( .B(arr[1005]), .A(arr[1046]), .S(n2982), .Y(n1668) );
  MUX2X1 U7234 ( .B(n1667), .A(n1664), .S(n3143), .Y(n1678) );
  MUX2X1 U7235 ( .B(arr[923]), .A(arr[964]), .S(n2982), .Y(n1672) );
  MUX2X1 U7236 ( .B(arr[841]), .A(arr[882]), .S(n2982), .Y(n1671) );
  MUX2X1 U7237 ( .B(arr[759]), .A(arr[800]), .S(n2982), .Y(n1675) );
  MUX2X1 U7238 ( .B(arr[677]), .A(arr[718]), .S(n2982), .Y(n1674) );
  MUX2X1 U7239 ( .B(n1673), .A(n1670), .S(n3143), .Y(n1677) );
  MUX2X1 U7240 ( .B(arr[595]), .A(arr[636]), .S(n2982), .Y(n1681) );
  MUX2X1 U7241 ( .B(arr[513]), .A(arr[554]), .S(n2982), .Y(n1680) );
  MUX2X1 U7242 ( .B(arr[431]), .A(arr[472]), .S(n2982), .Y(n1684) );
  MUX2X1 U7243 ( .B(arr[349]), .A(arr[390]), .S(n2982), .Y(n1683) );
  MUX2X1 U7244 ( .B(n1682), .A(n1679), .S(n3143), .Y(n1693) );
  MUX2X1 U7245 ( .B(arr[267]), .A(arr[308]), .S(n2983), .Y(n1687) );
  MUX2X1 U7246 ( .B(arr[185]), .A(arr[226]), .S(n2983), .Y(n1686) );
  MUX2X1 U7247 ( .B(arr[103]), .A(arr[144]), .S(n2983), .Y(n1690) );
  MUX2X1 U7248 ( .B(arr[21]), .A(arr[62]), .S(n2983), .Y(n1689) );
  MUX2X1 U7249 ( .B(n1688), .A(n1685), .S(n3143), .Y(n1692) );
  MUX2X1 U7250 ( .B(n1691), .A(n1676), .S(n3183), .Y(n1694) );
  MUX2X1 U7251 ( .B(arr[2564]), .A(arr[2605]), .S(n2983), .Y(n1698) );
  MUX2X1 U7252 ( .B(arr[2482]), .A(arr[2523]), .S(n2983), .Y(n1697) );
  MUX2X1 U7253 ( .B(arr[2400]), .A(arr[2441]), .S(n2983), .Y(n1701) );
  MUX2X1 U7254 ( .B(arr[2318]), .A(arr[2359]), .S(n2983), .Y(n1700) );
  MUX2X1 U7255 ( .B(n1699), .A(n1696), .S(n3143), .Y(n1710) );
  MUX2X1 U7256 ( .B(arr[2236]), .A(arr[2277]), .S(n2983), .Y(n1704) );
  MUX2X1 U7257 ( .B(arr[2154]), .A(arr[2195]), .S(n2983), .Y(n1703) );
  MUX2X1 U7258 ( .B(arr[2072]), .A(arr[2113]), .S(n2983), .Y(n1707) );
  MUX2X1 U7259 ( .B(arr[1990]), .A(arr[2031]), .S(n2983), .Y(n1706) );
  MUX2X1 U7260 ( .B(n1705), .A(n1702), .S(n3143), .Y(n1709) );
  MUX2X1 U7261 ( .B(arr[1908]), .A(arr[1949]), .S(n2984), .Y(n1713) );
  MUX2X1 U7262 ( .B(arr[1826]), .A(arr[1867]), .S(n2984), .Y(n1712) );
  MUX2X1 U7263 ( .B(arr[1744]), .A(arr[1785]), .S(n2984), .Y(n1716) );
  MUX2X1 U7264 ( .B(arr[1662]), .A(arr[1703]), .S(n2984), .Y(n1715) );
  MUX2X1 U7265 ( .B(n1714), .A(n1711), .S(n3143), .Y(n1725) );
  MUX2X1 U7266 ( .B(arr[1580]), .A(arr[1621]), .S(n2984), .Y(n1719) );
  MUX2X1 U7267 ( .B(arr[1498]), .A(arr[1539]), .S(n2984), .Y(n1718) );
  MUX2X1 U7268 ( .B(arr[1416]), .A(arr[1457]), .S(n2984), .Y(n1722) );
  MUX2X1 U7269 ( .B(arr[1334]), .A(arr[1375]), .S(n2984), .Y(n1721) );
  MUX2X1 U7270 ( .B(n1720), .A(n1717), .S(n3143), .Y(n1724) );
  MUX2X1 U7271 ( .B(n1723), .A(n1708), .S(n3183), .Y(n1757) );
  MUX2X1 U7272 ( .B(arr[1252]), .A(arr[1293]), .S(n2984), .Y(n1728) );
  MUX2X1 U7273 ( .B(arr[1170]), .A(arr[1211]), .S(n2984), .Y(n1727) );
  MUX2X1 U7274 ( .B(arr[1088]), .A(arr[1129]), .S(n2984), .Y(n1731) );
  MUX2X1 U7275 ( .B(arr[1006]), .A(arr[1047]), .S(n2984), .Y(n1730) );
  MUX2X1 U7276 ( .B(n1729), .A(n1726), .S(n3143), .Y(n1740) );
  MUX2X1 U7277 ( .B(arr[924]), .A(arr[965]), .S(n2985), .Y(n1734) );
  MUX2X1 U7278 ( .B(arr[842]), .A(arr[883]), .S(n2985), .Y(n1733) );
  MUX2X1 U7279 ( .B(arr[760]), .A(arr[801]), .S(n2985), .Y(n1737) );
  MUX2X1 U7280 ( .B(arr[678]), .A(arr[719]), .S(n2985), .Y(n1736) );
  MUX2X1 U7281 ( .B(n1735), .A(n1732), .S(n3143), .Y(n1739) );
  MUX2X1 U7282 ( .B(arr[596]), .A(arr[637]), .S(n2985), .Y(n1743) );
  MUX2X1 U7283 ( .B(arr[514]), .A(arr[555]), .S(n2985), .Y(n1742) );
  MUX2X1 U7284 ( .B(arr[432]), .A(arr[473]), .S(n2985), .Y(n1746) );
  MUX2X1 U7285 ( .B(arr[350]), .A(arr[391]), .S(n2985), .Y(n1745) );
  MUX2X1 U7286 ( .B(n1744), .A(n1741), .S(n3143), .Y(n1755) );
  MUX2X1 U7287 ( .B(arr[268]), .A(arr[309]), .S(n2985), .Y(n1749) );
  MUX2X1 U7288 ( .B(arr[186]), .A(arr[227]), .S(n2985), .Y(n1748) );
  MUX2X1 U7289 ( .B(arr[104]), .A(arr[145]), .S(n2985), .Y(n1752) );
  MUX2X1 U7290 ( .B(arr[22]), .A(arr[63]), .S(n2985), .Y(n1751) );
  MUX2X1 U7291 ( .B(n1750), .A(n1747), .S(n3143), .Y(n1754) );
  MUX2X1 U7292 ( .B(n1753), .A(n1738), .S(n3183), .Y(n1756) );
  MUX2X1 U7293 ( .B(arr[2565]), .A(arr[2606]), .S(n2986), .Y(n1760) );
  MUX2X1 U7294 ( .B(arr[2483]), .A(arr[2524]), .S(n2986), .Y(n1759) );
  MUX2X1 U7295 ( .B(arr[2401]), .A(arr[2442]), .S(n2986), .Y(n1763) );
  MUX2X1 U7296 ( .B(arr[2319]), .A(arr[2360]), .S(n2986), .Y(n1762) );
  MUX2X1 U7297 ( .B(n1761), .A(n1758), .S(n3144), .Y(n1772) );
  MUX2X1 U7298 ( .B(arr[2237]), .A(arr[2278]), .S(n2986), .Y(n1766) );
  MUX2X1 U7299 ( .B(arr[2155]), .A(arr[2196]), .S(n2986), .Y(n1765) );
  MUX2X1 U7300 ( .B(arr[2073]), .A(arr[2114]), .S(n2986), .Y(n1769) );
  MUX2X1 U7301 ( .B(arr[1991]), .A(arr[2032]), .S(n2986), .Y(n1768) );
  MUX2X1 U7302 ( .B(n1767), .A(n1764), .S(n3144), .Y(n1771) );
  MUX2X1 U7303 ( .B(arr[1909]), .A(arr[1950]), .S(n2986), .Y(n1775) );
  MUX2X1 U7304 ( .B(arr[1827]), .A(arr[1868]), .S(n2986), .Y(n1774) );
  MUX2X1 U7305 ( .B(arr[1745]), .A(arr[1786]), .S(n2986), .Y(n1778) );
  MUX2X1 U7306 ( .B(arr[1663]), .A(arr[1704]), .S(n2986), .Y(n1777) );
  MUX2X1 U7307 ( .B(n1776), .A(n1773), .S(n3144), .Y(n1787) );
  MUX2X1 U7308 ( .B(arr[1581]), .A(arr[1622]), .S(n2987), .Y(n1781) );
  MUX2X1 U7309 ( .B(arr[1499]), .A(arr[1540]), .S(n2987), .Y(n1780) );
  MUX2X1 U7310 ( .B(arr[1417]), .A(arr[1458]), .S(n2987), .Y(n1784) );
  MUX2X1 U7311 ( .B(arr[1335]), .A(arr[1376]), .S(n2987), .Y(n1783) );
  MUX2X1 U7312 ( .B(n1782), .A(n1779), .S(n3144), .Y(n1786) );
  MUX2X1 U7313 ( .B(n1785), .A(n1770), .S(n3184), .Y(n1819) );
  MUX2X1 U7314 ( .B(arr[1253]), .A(arr[1294]), .S(n2987), .Y(n1790) );
  MUX2X1 U7315 ( .B(arr[1171]), .A(arr[1212]), .S(n2987), .Y(n1789) );
  MUX2X1 U7316 ( .B(arr[1089]), .A(arr[1130]), .S(n2987), .Y(n1793) );
  MUX2X1 U7317 ( .B(arr[1007]), .A(arr[1048]), .S(n2987), .Y(n1792) );
  MUX2X1 U7318 ( .B(n1791), .A(n1788), .S(n3144), .Y(n1802) );
  MUX2X1 U7319 ( .B(arr[925]), .A(arr[966]), .S(n2987), .Y(n1796) );
  MUX2X1 U7320 ( .B(arr[843]), .A(arr[884]), .S(n2987), .Y(n1795) );
  MUX2X1 U7321 ( .B(arr[761]), .A(arr[802]), .S(n2987), .Y(n1799) );
  MUX2X1 U7322 ( .B(arr[679]), .A(arr[720]), .S(n2987), .Y(n1798) );
  MUX2X1 U7323 ( .B(n1797), .A(n1794), .S(n3144), .Y(n1801) );
  MUX2X1 U7324 ( .B(arr[597]), .A(arr[638]), .S(n2988), .Y(n1805) );
  MUX2X1 U7325 ( .B(arr[515]), .A(arr[556]), .S(n2988), .Y(n1804) );
  MUX2X1 U7326 ( .B(arr[433]), .A(arr[474]), .S(n2988), .Y(n1808) );
  MUX2X1 U7327 ( .B(arr[351]), .A(arr[392]), .S(n2988), .Y(n1807) );
  MUX2X1 U7328 ( .B(n1806), .A(n1803), .S(n3144), .Y(n1817) );
  MUX2X1 U7329 ( .B(arr[269]), .A(arr[310]), .S(n2988), .Y(n1811) );
  MUX2X1 U7330 ( .B(arr[187]), .A(arr[228]), .S(n2988), .Y(n1810) );
  MUX2X1 U7331 ( .B(arr[105]), .A(arr[146]), .S(n2988), .Y(n1814) );
  MUX2X1 U7332 ( .B(arr[23]), .A(arr[64]), .S(n2988), .Y(n1813) );
  MUX2X1 U7333 ( .B(n1812), .A(n1809), .S(n3144), .Y(n1816) );
  MUX2X1 U7334 ( .B(n1815), .A(n1800), .S(n3184), .Y(n1818) );
  MUX2X1 U7335 ( .B(arr[2566]), .A(arr[2607]), .S(n2988), .Y(n1822) );
  MUX2X1 U7336 ( .B(arr[2484]), .A(arr[2525]), .S(n2988), .Y(n1821) );
  MUX2X1 U7337 ( .B(arr[2402]), .A(arr[2443]), .S(n2988), .Y(n1825) );
  MUX2X1 U7338 ( .B(arr[2320]), .A(arr[2361]), .S(n2988), .Y(n1824) );
  MUX2X1 U7339 ( .B(n1823), .A(n1820), .S(n3144), .Y(n1834) );
  MUX2X1 U7340 ( .B(arr[2238]), .A(arr[2279]), .S(n2989), .Y(n1828) );
  MUX2X1 U7341 ( .B(arr[2156]), .A(arr[2197]), .S(n2989), .Y(n1827) );
  MUX2X1 U7342 ( .B(arr[2074]), .A(arr[2115]), .S(n2989), .Y(n1831) );
  MUX2X1 U7343 ( .B(arr[1992]), .A(arr[2033]), .S(n2989), .Y(n1830) );
  MUX2X1 U7344 ( .B(n1829), .A(n1826), .S(n3144), .Y(n1833) );
  MUX2X1 U7345 ( .B(arr[1910]), .A(arr[1951]), .S(n2989), .Y(n1837) );
  MUX2X1 U7346 ( .B(arr[1828]), .A(arr[1869]), .S(n2989), .Y(n1836) );
  MUX2X1 U7347 ( .B(arr[1746]), .A(arr[1787]), .S(n2989), .Y(n1840) );
  MUX2X1 U7348 ( .B(arr[1664]), .A(arr[1705]), .S(n2989), .Y(n1839) );
  MUX2X1 U7349 ( .B(n1838), .A(n1835), .S(n3144), .Y(n1849) );
  MUX2X1 U7350 ( .B(arr[1582]), .A(arr[1623]), .S(n2989), .Y(n1843) );
  MUX2X1 U7351 ( .B(arr[1500]), .A(arr[1541]), .S(n2989), .Y(n1842) );
  MUX2X1 U7352 ( .B(arr[1418]), .A(arr[1459]), .S(n2989), .Y(n1846) );
  MUX2X1 U7353 ( .B(arr[1336]), .A(arr[1377]), .S(n2989), .Y(n1845) );
  MUX2X1 U7354 ( .B(n1844), .A(n1841), .S(n3144), .Y(n1848) );
  MUX2X1 U7355 ( .B(n1847), .A(n1832), .S(n3184), .Y(n1881) );
  MUX2X1 U7356 ( .B(arr[1254]), .A(arr[1295]), .S(n2990), .Y(n1852) );
  MUX2X1 U7357 ( .B(arr[1172]), .A(arr[1213]), .S(n2990), .Y(n1851) );
  MUX2X1 U7358 ( .B(arr[1090]), .A(arr[1131]), .S(n2990), .Y(n1855) );
  MUX2X1 U7359 ( .B(arr[1008]), .A(arr[1049]), .S(n2990), .Y(n1854) );
  MUX2X1 U7360 ( .B(n1853), .A(n1850), .S(n3145), .Y(n1864) );
  MUX2X1 U7361 ( .B(arr[926]), .A(arr[967]), .S(n2990), .Y(n1858) );
  MUX2X1 U7362 ( .B(arr[844]), .A(arr[885]), .S(n2990), .Y(n1857) );
  MUX2X1 U7363 ( .B(arr[762]), .A(arr[803]), .S(n2990), .Y(n1861) );
  MUX2X1 U7364 ( .B(arr[680]), .A(arr[721]), .S(n2990), .Y(n1860) );
  MUX2X1 U7365 ( .B(n1859), .A(n1856), .S(n3145), .Y(n1863) );
  MUX2X1 U7366 ( .B(arr[598]), .A(arr[639]), .S(n2990), .Y(n1867) );
  MUX2X1 U7367 ( .B(arr[516]), .A(arr[557]), .S(n2990), .Y(n1866) );
  MUX2X1 U7368 ( .B(arr[434]), .A(arr[475]), .S(n2990), .Y(n1870) );
  MUX2X1 U7369 ( .B(arr[352]), .A(arr[393]), .S(n2990), .Y(n1869) );
  MUX2X1 U7370 ( .B(n1868), .A(n1865), .S(n3145), .Y(n1879) );
  MUX2X1 U7371 ( .B(arr[270]), .A(arr[311]), .S(n2991), .Y(n1873) );
  MUX2X1 U7372 ( .B(arr[188]), .A(arr[229]), .S(n2991), .Y(n1872) );
  MUX2X1 U7373 ( .B(arr[106]), .A(arr[147]), .S(n2991), .Y(n1876) );
  MUX2X1 U7374 ( .B(arr[24]), .A(arr[65]), .S(n2991), .Y(n1875) );
  MUX2X1 U7375 ( .B(n1874), .A(n1871), .S(n3145), .Y(n1878) );
  MUX2X1 U7376 ( .B(n1877), .A(n1862), .S(n3184), .Y(n1880) );
  MUX2X1 U7377 ( .B(arr[2567]), .A(arr[2608]), .S(n2991), .Y(n1884) );
  MUX2X1 U7378 ( .B(arr[2485]), .A(arr[2526]), .S(n2991), .Y(n1883) );
  MUX2X1 U7379 ( .B(arr[2403]), .A(arr[2444]), .S(n2991), .Y(n1887) );
  MUX2X1 U7380 ( .B(arr[2321]), .A(arr[2362]), .S(n2991), .Y(n1886) );
  MUX2X1 U7381 ( .B(n1885), .A(n1882), .S(n3145), .Y(n1896) );
  MUX2X1 U7382 ( .B(arr[2239]), .A(arr[2280]), .S(n2991), .Y(n1890) );
  MUX2X1 U7383 ( .B(arr[2157]), .A(arr[2198]), .S(n2991), .Y(n1889) );
  MUX2X1 U7384 ( .B(arr[2075]), .A(arr[2116]), .S(n2991), .Y(n1893) );
  MUX2X1 U7385 ( .B(arr[1993]), .A(arr[2034]), .S(n2991), .Y(n1892) );
  MUX2X1 U7386 ( .B(n1891), .A(n1888), .S(n3145), .Y(n1895) );
  MUX2X1 U7387 ( .B(arr[1911]), .A(arr[1952]), .S(n2992), .Y(n1899) );
  MUX2X1 U7388 ( .B(arr[1829]), .A(arr[1870]), .S(n2992), .Y(n1898) );
  MUX2X1 U7389 ( .B(arr[1747]), .A(arr[1788]), .S(n2992), .Y(n1902) );
  MUX2X1 U7390 ( .B(arr[1665]), .A(arr[1706]), .S(n2992), .Y(n1901) );
  MUX2X1 U7391 ( .B(n1900), .A(n1897), .S(n3145), .Y(n1911) );
  MUX2X1 U7392 ( .B(arr[1583]), .A(arr[1624]), .S(n2992), .Y(n1905) );
  MUX2X1 U7393 ( .B(arr[1501]), .A(arr[1542]), .S(n2992), .Y(n1904) );
  MUX2X1 U7394 ( .B(arr[1419]), .A(arr[1460]), .S(n2992), .Y(n1908) );
  MUX2X1 U7395 ( .B(arr[1337]), .A(arr[1378]), .S(n2992), .Y(n1907) );
  MUX2X1 U7396 ( .B(n1906), .A(n1903), .S(n3145), .Y(n1910) );
  MUX2X1 U7397 ( .B(n1909), .A(n1894), .S(n3184), .Y(n1943) );
  MUX2X1 U7398 ( .B(arr[1255]), .A(arr[1296]), .S(n2992), .Y(n1914) );
  MUX2X1 U7399 ( .B(arr[1173]), .A(arr[1214]), .S(n2992), .Y(n1913) );
  MUX2X1 U7400 ( .B(arr[1091]), .A(arr[1132]), .S(n2992), .Y(n1917) );
  MUX2X1 U7401 ( .B(arr[1009]), .A(arr[1050]), .S(n2992), .Y(n1916) );
  MUX2X1 U7402 ( .B(n1915), .A(n1912), .S(n3145), .Y(n1926) );
  MUX2X1 U7403 ( .B(arr[927]), .A(arr[968]), .S(n2993), .Y(n1920) );
  MUX2X1 U7404 ( .B(arr[845]), .A(arr[886]), .S(n2993), .Y(n1919) );
  MUX2X1 U7405 ( .B(arr[763]), .A(arr[804]), .S(n2993), .Y(n1923) );
  MUX2X1 U7406 ( .B(arr[681]), .A(arr[722]), .S(n2993), .Y(n1922) );
  MUX2X1 U7407 ( .B(n1921), .A(n1918), .S(n3145), .Y(n1925) );
  MUX2X1 U7408 ( .B(arr[599]), .A(arr[640]), .S(n2993), .Y(n1929) );
  MUX2X1 U7409 ( .B(arr[517]), .A(arr[558]), .S(n2993), .Y(n1928) );
  MUX2X1 U7410 ( .B(arr[435]), .A(arr[476]), .S(n2993), .Y(n1932) );
  MUX2X1 U7411 ( .B(arr[353]), .A(arr[394]), .S(n2993), .Y(n1931) );
  MUX2X1 U7412 ( .B(n1930), .A(n1927), .S(n3145), .Y(n1941) );
  MUX2X1 U7413 ( .B(arr[271]), .A(arr[312]), .S(n2993), .Y(n1935) );
  MUX2X1 U7414 ( .B(arr[189]), .A(arr[230]), .S(n2993), .Y(n1934) );
  MUX2X1 U7415 ( .B(arr[107]), .A(arr[148]), .S(n2993), .Y(n1938) );
  MUX2X1 U7416 ( .B(arr[25]), .A(arr[66]), .S(n2993), .Y(n1937) );
  MUX2X1 U7417 ( .B(n1936), .A(n1933), .S(n3145), .Y(n1940) );
  MUX2X1 U7418 ( .B(n1939), .A(n1924), .S(n3184), .Y(n1942) );
  MUX2X1 U7419 ( .B(arr[2568]), .A(arr[2609]), .S(n2994), .Y(n1946) );
  MUX2X1 U7420 ( .B(arr[2486]), .A(arr[2527]), .S(n2994), .Y(n1945) );
  MUX2X1 U7421 ( .B(arr[2404]), .A(arr[2445]), .S(n2994), .Y(n1949) );
  MUX2X1 U7422 ( .B(arr[2322]), .A(arr[2363]), .S(n2994), .Y(n1948) );
  MUX2X1 U7423 ( .B(n1947), .A(n1944), .S(n3146), .Y(n1958) );
  MUX2X1 U7424 ( .B(arr[2240]), .A(arr[2281]), .S(n2994), .Y(n1952) );
  MUX2X1 U7425 ( .B(arr[2158]), .A(arr[2199]), .S(n2994), .Y(n1951) );
  MUX2X1 U7426 ( .B(arr[2076]), .A(arr[2117]), .S(n2994), .Y(n1955) );
  MUX2X1 U7427 ( .B(arr[1994]), .A(arr[2035]), .S(n2994), .Y(n1954) );
  MUX2X1 U7428 ( .B(n1953), .A(n1950), .S(n3146), .Y(n1957) );
  MUX2X1 U7429 ( .B(arr[1912]), .A(arr[1953]), .S(n2994), .Y(n1961) );
  MUX2X1 U7430 ( .B(arr[1830]), .A(arr[1871]), .S(n2994), .Y(n1960) );
  MUX2X1 U7431 ( .B(arr[1748]), .A(arr[1789]), .S(n2994), .Y(n1964) );
  MUX2X1 U7432 ( .B(arr[1666]), .A(arr[1707]), .S(n2994), .Y(n1963) );
  MUX2X1 U7433 ( .B(n1962), .A(n1959), .S(n3146), .Y(n1973) );
  MUX2X1 U7434 ( .B(arr[1584]), .A(arr[1625]), .S(n2995), .Y(n1967) );
  MUX2X1 U7435 ( .B(arr[1502]), .A(arr[1543]), .S(n2995), .Y(n1966) );
  MUX2X1 U7436 ( .B(arr[1420]), .A(arr[1461]), .S(n2995), .Y(n1970) );
  MUX2X1 U7437 ( .B(arr[1338]), .A(arr[1379]), .S(n2995), .Y(n1969) );
  MUX2X1 U7438 ( .B(n1968), .A(n1965), .S(n3146), .Y(n1972) );
  MUX2X1 U7439 ( .B(n1971), .A(n1956), .S(n3184), .Y(n2005) );
  MUX2X1 U7440 ( .B(arr[1256]), .A(arr[1297]), .S(n2995), .Y(n1976) );
  MUX2X1 U7441 ( .B(arr[1174]), .A(arr[1215]), .S(n2995), .Y(n1975) );
  MUX2X1 U7442 ( .B(arr[1092]), .A(arr[1133]), .S(n2995), .Y(n1979) );
  MUX2X1 U7443 ( .B(arr[1010]), .A(arr[1051]), .S(n2995), .Y(n1978) );
  MUX2X1 U7444 ( .B(n1977), .A(n1974), .S(n3146), .Y(n1988) );
  MUX2X1 U7445 ( .B(arr[928]), .A(arr[969]), .S(n2995), .Y(n1982) );
  MUX2X1 U7446 ( .B(arr[846]), .A(arr[887]), .S(n2995), .Y(n1981) );
  MUX2X1 U7447 ( .B(arr[764]), .A(arr[805]), .S(n2995), .Y(n1985) );
  MUX2X1 U7448 ( .B(arr[682]), .A(arr[723]), .S(n2995), .Y(n1984) );
  MUX2X1 U7449 ( .B(n1983), .A(n1980), .S(n3146), .Y(n1987) );
  MUX2X1 U7450 ( .B(arr[600]), .A(arr[641]), .S(n2996), .Y(n1991) );
  MUX2X1 U7451 ( .B(arr[518]), .A(arr[559]), .S(n2996), .Y(n1990) );
  MUX2X1 U7452 ( .B(arr[436]), .A(arr[477]), .S(n2996), .Y(n1994) );
  MUX2X1 U7453 ( .B(arr[354]), .A(arr[395]), .S(n2996), .Y(n1993) );
  MUX2X1 U7454 ( .B(n1992), .A(n1989), .S(n3146), .Y(n2003) );
  MUX2X1 U7455 ( .B(arr[272]), .A(arr[313]), .S(n2996), .Y(n1997) );
  MUX2X1 U7456 ( .B(arr[190]), .A(arr[231]), .S(n2996), .Y(n1996) );
  MUX2X1 U7457 ( .B(arr[108]), .A(arr[149]), .S(n2996), .Y(n2000) );
  MUX2X1 U7458 ( .B(arr[26]), .A(arr[67]), .S(n2996), .Y(n1999) );
  MUX2X1 U7459 ( .B(n1998), .A(n1995), .S(n3146), .Y(n2002) );
  MUX2X1 U7460 ( .B(n2001), .A(n1986), .S(n3184), .Y(n2004) );
  MUX2X1 U7461 ( .B(arr[2569]), .A(arr[2610]), .S(n2996), .Y(n2008) );
  MUX2X1 U7462 ( .B(arr[2487]), .A(arr[2528]), .S(n2996), .Y(n2007) );
  MUX2X1 U7463 ( .B(arr[2405]), .A(arr[2446]), .S(n2996), .Y(n2011) );
  MUX2X1 U7464 ( .B(arr[2323]), .A(arr[2364]), .S(n2996), .Y(n2010) );
  MUX2X1 U7465 ( .B(n2009), .A(n2006), .S(n3146), .Y(n2020) );
  MUX2X1 U7466 ( .B(arr[2241]), .A(arr[2282]), .S(n2997), .Y(n2014) );
  MUX2X1 U7467 ( .B(arr[2159]), .A(arr[2200]), .S(n2997), .Y(n2013) );
  MUX2X1 U7468 ( .B(arr[2077]), .A(arr[2118]), .S(n2997), .Y(n2017) );
  MUX2X1 U7469 ( .B(arr[1995]), .A(arr[2036]), .S(n2997), .Y(n2016) );
  MUX2X1 U7470 ( .B(n2015), .A(n2012), .S(n3146), .Y(n2019) );
  MUX2X1 U7471 ( .B(arr[1913]), .A(arr[1954]), .S(n2997), .Y(n2023) );
  MUX2X1 U7472 ( .B(arr[1831]), .A(arr[1872]), .S(n2997), .Y(n2022) );
  MUX2X1 U7473 ( .B(arr[1749]), .A(arr[1790]), .S(n2997), .Y(n2026) );
  MUX2X1 U7474 ( .B(arr[1667]), .A(arr[1708]), .S(n2997), .Y(n2025) );
  MUX2X1 U7475 ( .B(n2024), .A(n2021), .S(n3146), .Y(n2035) );
  MUX2X1 U7476 ( .B(arr[1585]), .A(arr[1626]), .S(n2997), .Y(n2029) );
  MUX2X1 U7477 ( .B(arr[1503]), .A(arr[1544]), .S(n2997), .Y(n2028) );
  MUX2X1 U7478 ( .B(arr[1421]), .A(arr[1462]), .S(n2997), .Y(n2032) );
  MUX2X1 U7479 ( .B(arr[1339]), .A(arr[1380]), .S(n2997), .Y(n2031) );
  MUX2X1 U7480 ( .B(n2030), .A(n2027), .S(n3146), .Y(n2034) );
  MUX2X1 U7481 ( .B(n2033), .A(n2018), .S(n3184), .Y(n2067) );
  MUX2X1 U7482 ( .B(arr[1257]), .A(arr[1298]), .S(n2998), .Y(n2038) );
  MUX2X1 U7483 ( .B(arr[1175]), .A(arr[1216]), .S(n2998), .Y(n2037) );
  MUX2X1 U7484 ( .B(arr[1093]), .A(arr[1134]), .S(n2998), .Y(n2041) );
  MUX2X1 U7485 ( .B(arr[1011]), .A(arr[1052]), .S(n2998), .Y(n2040) );
  MUX2X1 U7486 ( .B(n2039), .A(n2036), .S(n3147), .Y(n2050) );
  MUX2X1 U7487 ( .B(arr[929]), .A(arr[970]), .S(n2998), .Y(n2044) );
  MUX2X1 U7488 ( .B(arr[847]), .A(arr[888]), .S(n2998), .Y(n2043) );
  MUX2X1 U7489 ( .B(arr[765]), .A(arr[806]), .S(n2998), .Y(n2047) );
  MUX2X1 U7490 ( .B(arr[683]), .A(arr[724]), .S(n2998), .Y(n2046) );
  MUX2X1 U7491 ( .B(n2045), .A(n2042), .S(n3147), .Y(n2049) );
  MUX2X1 U7492 ( .B(arr[601]), .A(arr[642]), .S(n2998), .Y(n2053) );
  MUX2X1 U7493 ( .B(arr[519]), .A(arr[560]), .S(n2998), .Y(n2052) );
  MUX2X1 U7494 ( .B(arr[437]), .A(arr[478]), .S(n2998), .Y(n2056) );
  MUX2X1 U7495 ( .B(arr[355]), .A(arr[396]), .S(n2998), .Y(n2055) );
  MUX2X1 U7496 ( .B(n2054), .A(n2051), .S(n3147), .Y(n2065) );
  MUX2X1 U7497 ( .B(arr[273]), .A(arr[314]), .S(n2999), .Y(n2059) );
  MUX2X1 U7498 ( .B(arr[191]), .A(arr[232]), .S(n2999), .Y(n2058) );
  MUX2X1 U7499 ( .B(arr[109]), .A(arr[150]), .S(n2999), .Y(n2062) );
  MUX2X1 U7500 ( .B(arr[27]), .A(arr[68]), .S(n2999), .Y(n2061) );
  MUX2X1 U7501 ( .B(n2060), .A(n2057), .S(n3147), .Y(n2064) );
  MUX2X1 U7502 ( .B(n2063), .A(n2048), .S(n3184), .Y(n2066) );
  MUX2X1 U7503 ( .B(arr[2570]), .A(arr[2611]), .S(n2999), .Y(n2070) );
  MUX2X1 U7504 ( .B(arr[2488]), .A(arr[2529]), .S(n2999), .Y(n2069) );
  MUX2X1 U7505 ( .B(arr[2406]), .A(arr[2447]), .S(n2999), .Y(n2073) );
  MUX2X1 U7506 ( .B(arr[2324]), .A(arr[2365]), .S(n2999), .Y(n2072) );
  MUX2X1 U7507 ( .B(n2071), .A(n2068), .S(n3147), .Y(n2082) );
  MUX2X1 U7508 ( .B(arr[2242]), .A(arr[2283]), .S(n2999), .Y(n2076) );
  MUX2X1 U7509 ( .B(arr[2160]), .A(arr[2201]), .S(n2999), .Y(n2075) );
  MUX2X1 U7510 ( .B(arr[2078]), .A(arr[2119]), .S(n2999), .Y(n2079) );
  MUX2X1 U7511 ( .B(arr[1996]), .A(arr[2037]), .S(n2999), .Y(n2078) );
  MUX2X1 U7512 ( .B(n2077), .A(n2074), .S(n3147), .Y(n2081) );
  MUX2X1 U7513 ( .B(arr[1914]), .A(arr[1955]), .S(n3000), .Y(n2085) );
  MUX2X1 U7514 ( .B(arr[1832]), .A(arr[1873]), .S(n3000), .Y(n2084) );
  MUX2X1 U7515 ( .B(arr[1750]), .A(arr[1791]), .S(n3000), .Y(n2088) );
  MUX2X1 U7516 ( .B(arr[1668]), .A(arr[1709]), .S(n3000), .Y(n2087) );
  MUX2X1 U7517 ( .B(n2086), .A(n2083), .S(n3147), .Y(n2097) );
  MUX2X1 U7518 ( .B(arr[1586]), .A(arr[1627]), .S(n3000), .Y(n2091) );
  MUX2X1 U7519 ( .B(arr[1504]), .A(arr[1545]), .S(n3000), .Y(n2090) );
  MUX2X1 U7520 ( .B(arr[1422]), .A(arr[1463]), .S(n3000), .Y(n2094) );
  MUX2X1 U7521 ( .B(arr[1340]), .A(arr[1381]), .S(n3000), .Y(n2093) );
  MUX2X1 U7522 ( .B(n2092), .A(n2089), .S(n3147), .Y(n2096) );
  MUX2X1 U7523 ( .B(n2095), .A(n2080), .S(n3184), .Y(n2129) );
  MUX2X1 U7524 ( .B(arr[1258]), .A(arr[1299]), .S(n3000), .Y(n2100) );
  MUX2X1 U7525 ( .B(arr[1176]), .A(arr[1217]), .S(n3000), .Y(n2099) );
  MUX2X1 U7526 ( .B(arr[1094]), .A(arr[1135]), .S(n3000), .Y(n2103) );
  MUX2X1 U7527 ( .B(arr[1012]), .A(arr[1053]), .S(n3000), .Y(n2102) );
  MUX2X1 U7528 ( .B(n2101), .A(n2098), .S(n3147), .Y(n2112) );
  MUX2X1 U7529 ( .B(arr[930]), .A(arr[971]), .S(n3001), .Y(n2106) );
  MUX2X1 U7530 ( .B(arr[848]), .A(arr[889]), .S(n3001), .Y(n2105) );
  MUX2X1 U7531 ( .B(arr[766]), .A(arr[807]), .S(n3001), .Y(n2109) );
  MUX2X1 U7532 ( .B(arr[684]), .A(arr[725]), .S(n3001), .Y(n2108) );
  MUX2X1 U7533 ( .B(n2107), .A(n2104), .S(n3147), .Y(n2111) );
  MUX2X1 U7534 ( .B(arr[602]), .A(arr[643]), .S(n3001), .Y(n2115) );
  MUX2X1 U7535 ( .B(arr[520]), .A(arr[561]), .S(n3001), .Y(n2114) );
  MUX2X1 U7536 ( .B(arr[438]), .A(arr[479]), .S(n3001), .Y(n2118) );
  MUX2X1 U7537 ( .B(arr[356]), .A(arr[397]), .S(n3001), .Y(n2117) );
  MUX2X1 U7538 ( .B(n2116), .A(n2113), .S(n3147), .Y(n2127) );
  MUX2X1 U7539 ( .B(arr[274]), .A(arr[315]), .S(n3001), .Y(n2121) );
  MUX2X1 U7540 ( .B(arr[192]), .A(arr[233]), .S(n3001), .Y(n2120) );
  MUX2X1 U7541 ( .B(arr[110]), .A(arr[151]), .S(n3001), .Y(n2124) );
  MUX2X1 U7542 ( .B(arr[28]), .A(arr[69]), .S(n3001), .Y(n2123) );
  MUX2X1 U7543 ( .B(n2122), .A(n2119), .S(n3147), .Y(n2126) );
  MUX2X1 U7544 ( .B(n2125), .A(n2110), .S(n3184), .Y(n2128) );
  MUX2X1 U7545 ( .B(arr[2571]), .A(arr[2612]), .S(n3002), .Y(n2132) );
  MUX2X1 U7546 ( .B(arr[2489]), .A(arr[2530]), .S(n3002), .Y(n2131) );
  MUX2X1 U7547 ( .B(arr[2407]), .A(arr[2448]), .S(n3002), .Y(n2135) );
  MUX2X1 U7548 ( .B(arr[2325]), .A(arr[2366]), .S(n3002), .Y(n2134) );
  MUX2X1 U7549 ( .B(n2133), .A(n2130), .S(n3148), .Y(n2144) );
  MUX2X1 U7550 ( .B(arr[2243]), .A(arr[2284]), .S(n3002), .Y(n2138) );
  MUX2X1 U7551 ( .B(arr[2161]), .A(arr[2202]), .S(n3002), .Y(n2137) );
  MUX2X1 U7552 ( .B(arr[2079]), .A(arr[2120]), .S(n3002), .Y(n2141) );
  MUX2X1 U7553 ( .B(arr[1997]), .A(arr[2038]), .S(n3002), .Y(n2140) );
  MUX2X1 U7554 ( .B(n2139), .A(n2136), .S(n3148), .Y(n2143) );
  MUX2X1 U7555 ( .B(arr[1915]), .A(arr[1956]), .S(n3002), .Y(n2147) );
  MUX2X1 U7556 ( .B(arr[1833]), .A(arr[1874]), .S(n3002), .Y(n2146) );
  MUX2X1 U7557 ( .B(arr[1751]), .A(arr[1792]), .S(n3002), .Y(n2150) );
  MUX2X1 U7558 ( .B(arr[1669]), .A(arr[1710]), .S(n3002), .Y(n2149) );
  MUX2X1 U7559 ( .B(n2148), .A(n2145), .S(n3148), .Y(n2159) );
  MUX2X1 U7560 ( .B(arr[1587]), .A(arr[1628]), .S(n3003), .Y(n2153) );
  MUX2X1 U7561 ( .B(arr[1505]), .A(arr[1546]), .S(n3003), .Y(n2152) );
  MUX2X1 U7562 ( .B(arr[1423]), .A(arr[1464]), .S(n3003), .Y(n2156) );
  MUX2X1 U7563 ( .B(arr[1341]), .A(arr[1382]), .S(n3003), .Y(n2155) );
  MUX2X1 U7564 ( .B(n2154), .A(n2151), .S(n3148), .Y(n2158) );
  MUX2X1 U7565 ( .B(n2157), .A(n2142), .S(n3185), .Y(n2191) );
  MUX2X1 U7566 ( .B(arr[1259]), .A(arr[1300]), .S(n3003), .Y(n2162) );
  MUX2X1 U7567 ( .B(arr[1177]), .A(arr[1218]), .S(n3003), .Y(n2161) );
  MUX2X1 U7568 ( .B(arr[1095]), .A(arr[1136]), .S(n3003), .Y(n2165) );
  MUX2X1 U7569 ( .B(arr[1013]), .A(arr[1054]), .S(n3003), .Y(n2164) );
  MUX2X1 U7570 ( .B(n2163), .A(n2160), .S(n3148), .Y(n2174) );
  MUX2X1 U7571 ( .B(arr[931]), .A(arr[972]), .S(n3003), .Y(n2168) );
  MUX2X1 U7572 ( .B(arr[849]), .A(arr[890]), .S(n3003), .Y(n2167) );
  MUX2X1 U7573 ( .B(arr[767]), .A(arr[808]), .S(n3003), .Y(n2171) );
  MUX2X1 U7574 ( .B(arr[685]), .A(arr[726]), .S(n3003), .Y(n2170) );
  MUX2X1 U7575 ( .B(n2169), .A(n2166), .S(n3148), .Y(n2173) );
  MUX2X1 U7576 ( .B(arr[603]), .A(arr[644]), .S(n3004), .Y(n2177) );
  MUX2X1 U7577 ( .B(arr[521]), .A(arr[562]), .S(n3004), .Y(n2176) );
  MUX2X1 U7578 ( .B(arr[439]), .A(arr[480]), .S(n3004), .Y(n2180) );
  MUX2X1 U7579 ( .B(arr[357]), .A(arr[398]), .S(n3004), .Y(n2179) );
  MUX2X1 U7580 ( .B(n2178), .A(n2175), .S(n3148), .Y(n2189) );
  MUX2X1 U7581 ( .B(arr[275]), .A(arr[316]), .S(n3004), .Y(n2183) );
  MUX2X1 U7582 ( .B(arr[193]), .A(arr[234]), .S(n3004), .Y(n2182) );
  MUX2X1 U7583 ( .B(arr[111]), .A(arr[152]), .S(n3004), .Y(n2186) );
  MUX2X1 U7584 ( .B(arr[29]), .A(arr[70]), .S(n3004), .Y(n2185) );
  MUX2X1 U7585 ( .B(n2184), .A(n2181), .S(n3148), .Y(n2188) );
  MUX2X1 U7586 ( .B(n2187), .A(n2172), .S(n3185), .Y(n2190) );
  MUX2X1 U7587 ( .B(arr[2572]), .A(arr[2613]), .S(n3004), .Y(n2194) );
  MUX2X1 U7588 ( .B(arr[2490]), .A(arr[2531]), .S(n3004), .Y(n2193) );
  MUX2X1 U7589 ( .B(arr[2408]), .A(arr[2449]), .S(n3004), .Y(n2197) );
  MUX2X1 U7590 ( .B(arr[2326]), .A(arr[2367]), .S(n3004), .Y(n2196) );
  MUX2X1 U7591 ( .B(n2195), .A(n2192), .S(n3148), .Y(n2206) );
  MUX2X1 U7592 ( .B(arr[2244]), .A(arr[2285]), .S(n3005), .Y(n2200) );
  MUX2X1 U7593 ( .B(arr[2162]), .A(arr[2203]), .S(n3005), .Y(n2199) );
  MUX2X1 U7594 ( .B(arr[2080]), .A(arr[2121]), .S(n3005), .Y(n2203) );
  MUX2X1 U7595 ( .B(arr[1998]), .A(arr[2039]), .S(n3005), .Y(n2202) );
  MUX2X1 U7596 ( .B(n2201), .A(n2198), .S(n3148), .Y(n2205) );
  MUX2X1 U7597 ( .B(arr[1916]), .A(arr[1957]), .S(n3005), .Y(n2209) );
  MUX2X1 U7598 ( .B(arr[1834]), .A(arr[1875]), .S(n3005), .Y(n2208) );
  MUX2X1 U7599 ( .B(arr[1752]), .A(arr[1793]), .S(n3005), .Y(n2212) );
  MUX2X1 U7600 ( .B(arr[1670]), .A(arr[1711]), .S(n3005), .Y(n2211) );
  MUX2X1 U7601 ( .B(n2210), .A(n2207), .S(n3148), .Y(n2221) );
  MUX2X1 U7602 ( .B(arr[1588]), .A(arr[1629]), .S(n3005), .Y(n2215) );
  MUX2X1 U7603 ( .B(arr[1506]), .A(arr[1547]), .S(n3005), .Y(n2214) );
  MUX2X1 U7604 ( .B(arr[1424]), .A(arr[1465]), .S(n3005), .Y(n2218) );
  MUX2X1 U7605 ( .B(arr[1342]), .A(arr[1383]), .S(n3005), .Y(n2217) );
  MUX2X1 U7606 ( .B(n2216), .A(n2213), .S(n3148), .Y(n2220) );
  MUX2X1 U7607 ( .B(n2219), .A(n2204), .S(n3185), .Y(n2253) );
  MUX2X1 U7608 ( .B(arr[1260]), .A(arr[1301]), .S(n3006), .Y(n2224) );
  MUX2X1 U7609 ( .B(arr[1178]), .A(arr[1219]), .S(n3006), .Y(n2223) );
  MUX2X1 U7610 ( .B(arr[1096]), .A(arr[1137]), .S(n3006), .Y(n2227) );
  MUX2X1 U7611 ( .B(arr[1014]), .A(arr[1055]), .S(n3006), .Y(n2226) );
  MUX2X1 U7612 ( .B(n2225), .A(n2222), .S(n3149), .Y(n2236) );
  MUX2X1 U7613 ( .B(arr[932]), .A(arr[973]), .S(n3006), .Y(n2230) );
  MUX2X1 U7614 ( .B(arr[850]), .A(arr[891]), .S(n3006), .Y(n2229) );
  MUX2X1 U7615 ( .B(arr[768]), .A(arr[809]), .S(n3006), .Y(n2233) );
  MUX2X1 U7616 ( .B(arr[686]), .A(arr[727]), .S(n3006), .Y(n2232) );
  MUX2X1 U7617 ( .B(n2231), .A(n2228), .S(n3149), .Y(n2235) );
  MUX2X1 U7618 ( .B(arr[604]), .A(arr[645]), .S(n3006), .Y(n2239) );
  MUX2X1 U7619 ( .B(arr[522]), .A(arr[563]), .S(n3006), .Y(n2238) );
  MUX2X1 U7620 ( .B(arr[440]), .A(arr[481]), .S(n3006), .Y(n2242) );
  MUX2X1 U7621 ( .B(arr[358]), .A(arr[399]), .S(n3006), .Y(n2241) );
  MUX2X1 U7622 ( .B(n2240), .A(n2237), .S(n3149), .Y(n2251) );
  MUX2X1 U7623 ( .B(arr[276]), .A(arr[317]), .S(n3007), .Y(n2245) );
  MUX2X1 U7624 ( .B(arr[194]), .A(arr[235]), .S(n3007), .Y(n2244) );
  MUX2X1 U7625 ( .B(arr[112]), .A(arr[153]), .S(n3007), .Y(n2248) );
  MUX2X1 U7626 ( .B(arr[30]), .A(arr[71]), .S(n3007), .Y(n2247) );
  MUX2X1 U7627 ( .B(n2246), .A(n2243), .S(n3149), .Y(n2250) );
  MUX2X1 U7628 ( .B(n2249), .A(n2234), .S(n3185), .Y(n2252) );
  MUX2X1 U7629 ( .B(arr[2573]), .A(arr[2614]), .S(n3007), .Y(n2256) );
  MUX2X1 U7630 ( .B(arr[2491]), .A(arr[2532]), .S(n3007), .Y(n2255) );
  MUX2X1 U7631 ( .B(arr[2409]), .A(arr[2450]), .S(n3007), .Y(n2259) );
  MUX2X1 U7632 ( .B(arr[2327]), .A(arr[2368]), .S(n3007), .Y(n2258) );
  MUX2X1 U7633 ( .B(n2257), .A(n2254), .S(n3149), .Y(n2268) );
  MUX2X1 U7634 ( .B(arr[2245]), .A(arr[2286]), .S(n3007), .Y(n2262) );
  MUX2X1 U7635 ( .B(arr[2163]), .A(arr[2204]), .S(n3007), .Y(n2261) );
  MUX2X1 U7636 ( .B(arr[2081]), .A(arr[2122]), .S(n3007), .Y(n2265) );
  MUX2X1 U7637 ( .B(arr[1999]), .A(arr[2040]), .S(n3007), .Y(n2264) );
  MUX2X1 U7638 ( .B(n2263), .A(n2260), .S(n3149), .Y(n2267) );
  MUX2X1 U7639 ( .B(arr[1917]), .A(arr[1958]), .S(n3008), .Y(n2271) );
  MUX2X1 U7640 ( .B(arr[1835]), .A(arr[1876]), .S(n3008), .Y(n2270) );
  MUX2X1 U7641 ( .B(arr[1753]), .A(arr[1794]), .S(n3008), .Y(n2274) );
  MUX2X1 U7642 ( .B(arr[1671]), .A(arr[1712]), .S(n3008), .Y(n2273) );
  MUX2X1 U7643 ( .B(n2272), .A(n2269), .S(n3149), .Y(n2283) );
  MUX2X1 U7644 ( .B(arr[1589]), .A(arr[1630]), .S(n3008), .Y(n2277) );
  MUX2X1 U7645 ( .B(arr[1507]), .A(arr[1548]), .S(n3008), .Y(n2276) );
  MUX2X1 U7646 ( .B(arr[1425]), .A(arr[1466]), .S(n3008), .Y(n2280) );
  MUX2X1 U7647 ( .B(arr[1343]), .A(arr[1384]), .S(n3008), .Y(n2279) );
  MUX2X1 U7648 ( .B(n2278), .A(n2275), .S(n3149), .Y(n2282) );
  MUX2X1 U7649 ( .B(n2281), .A(n2266), .S(n3185), .Y(n2315) );
  MUX2X1 U7650 ( .B(arr[1261]), .A(arr[1302]), .S(n3008), .Y(n2286) );
  MUX2X1 U7651 ( .B(arr[1179]), .A(arr[1220]), .S(n3008), .Y(n2285) );
  MUX2X1 U7652 ( .B(arr[1097]), .A(arr[1138]), .S(n3008), .Y(n2289) );
  MUX2X1 U7653 ( .B(arr[1015]), .A(arr[1056]), .S(n3008), .Y(n2288) );
  MUX2X1 U7654 ( .B(n2287), .A(n2284), .S(n3149), .Y(n2298) );
  MUX2X1 U7655 ( .B(arr[933]), .A(arr[974]), .S(n3009), .Y(n2292) );
  MUX2X1 U7656 ( .B(arr[851]), .A(arr[892]), .S(n3009), .Y(n2291) );
  MUX2X1 U7657 ( .B(arr[769]), .A(arr[810]), .S(n3009), .Y(n2295) );
  MUX2X1 U7658 ( .B(arr[687]), .A(arr[728]), .S(n3009), .Y(n2294) );
  MUX2X1 U7659 ( .B(n2293), .A(n2290), .S(n3149), .Y(n2297) );
  MUX2X1 U7660 ( .B(arr[605]), .A(arr[646]), .S(n3009), .Y(n2301) );
  MUX2X1 U7661 ( .B(arr[523]), .A(arr[564]), .S(n3009), .Y(n2300) );
  MUX2X1 U7662 ( .B(arr[441]), .A(arr[482]), .S(n3009), .Y(n2304) );
  MUX2X1 U7663 ( .B(arr[359]), .A(arr[400]), .S(n3009), .Y(n2303) );
  MUX2X1 U7664 ( .B(n2302), .A(n2299), .S(n3149), .Y(n2313) );
  MUX2X1 U7665 ( .B(arr[277]), .A(arr[318]), .S(n3009), .Y(n2307) );
  MUX2X1 U7666 ( .B(arr[195]), .A(arr[236]), .S(n3009), .Y(n2306) );
  MUX2X1 U7667 ( .B(arr[113]), .A(arr[154]), .S(n3009), .Y(n2310) );
  MUX2X1 U7668 ( .B(arr[31]), .A(arr[72]), .S(n3009), .Y(n2309) );
  MUX2X1 U7669 ( .B(n2308), .A(n2305), .S(n3149), .Y(n2312) );
  MUX2X1 U7670 ( .B(n2311), .A(n2296), .S(n3185), .Y(n2314) );
  MUX2X1 U7671 ( .B(arr[2574]), .A(arr[2615]), .S(n3010), .Y(n2318) );
  MUX2X1 U7672 ( .B(arr[2492]), .A(arr[2533]), .S(n3010), .Y(n2317) );
  MUX2X1 U7673 ( .B(arr[2410]), .A(arr[2451]), .S(n3010), .Y(n2321) );
  MUX2X1 U7674 ( .B(arr[2328]), .A(arr[2369]), .S(n3010), .Y(n2320) );
  MUX2X1 U7675 ( .B(n2319), .A(n2316), .S(n3150), .Y(n2330) );
  MUX2X1 U7676 ( .B(arr[2246]), .A(arr[2287]), .S(n3010), .Y(n2324) );
  MUX2X1 U7677 ( .B(arr[2164]), .A(arr[2205]), .S(n3010), .Y(n2323) );
  MUX2X1 U7678 ( .B(arr[2082]), .A(arr[2123]), .S(n3010), .Y(n2327) );
  MUX2X1 U7679 ( .B(arr[2000]), .A(arr[2041]), .S(n3010), .Y(n2326) );
  MUX2X1 U7680 ( .B(n2325), .A(n2322), .S(n3150), .Y(n2329) );
  MUX2X1 U7681 ( .B(arr[1918]), .A(arr[1959]), .S(n3010), .Y(n2333) );
  MUX2X1 U7682 ( .B(arr[1836]), .A(arr[1877]), .S(n3010), .Y(n2332) );
  MUX2X1 U7683 ( .B(arr[1754]), .A(arr[1795]), .S(n3010), .Y(n2336) );
  MUX2X1 U7684 ( .B(arr[1672]), .A(arr[1713]), .S(n3010), .Y(n2335) );
  MUX2X1 U7685 ( .B(n2334), .A(n2331), .S(n3150), .Y(n2345) );
  MUX2X1 U7686 ( .B(arr[1590]), .A(arr[1631]), .S(n3011), .Y(n2339) );
  MUX2X1 U7687 ( .B(arr[1508]), .A(arr[1549]), .S(n3011), .Y(n2338) );
  MUX2X1 U7688 ( .B(arr[1426]), .A(arr[1467]), .S(n3011), .Y(n2342) );
  MUX2X1 U7689 ( .B(arr[1344]), .A(arr[1385]), .S(n3011), .Y(n2341) );
  MUX2X1 U7690 ( .B(n2340), .A(n2337), .S(n3150), .Y(n2344) );
  MUX2X1 U7691 ( .B(n2343), .A(n2328), .S(n3185), .Y(n2377) );
  MUX2X1 U7692 ( .B(arr[1262]), .A(arr[1303]), .S(n3011), .Y(n2348) );
  MUX2X1 U7693 ( .B(arr[1180]), .A(arr[1221]), .S(n3011), .Y(n2347) );
  MUX2X1 U7694 ( .B(arr[1098]), .A(arr[1139]), .S(n3011), .Y(n2351) );
  MUX2X1 U7695 ( .B(arr[1016]), .A(arr[1057]), .S(n3011), .Y(n2350) );
  MUX2X1 U7696 ( .B(n2349), .A(n2346), .S(n3150), .Y(n2360) );
  MUX2X1 U7697 ( .B(arr[934]), .A(arr[975]), .S(n3011), .Y(n2354) );
  MUX2X1 U7698 ( .B(arr[852]), .A(arr[893]), .S(n3011), .Y(n2353) );
  MUX2X1 U7699 ( .B(arr[770]), .A(arr[811]), .S(n3011), .Y(n2357) );
  MUX2X1 U7700 ( .B(arr[688]), .A(arr[729]), .S(n3011), .Y(n2356) );
  MUX2X1 U7701 ( .B(n2355), .A(n2352), .S(n3150), .Y(n2359) );
  MUX2X1 U7702 ( .B(arr[606]), .A(arr[647]), .S(n3012), .Y(n2363) );
  MUX2X1 U7703 ( .B(arr[524]), .A(arr[565]), .S(n3012), .Y(n2362) );
  MUX2X1 U7704 ( .B(arr[442]), .A(arr[483]), .S(n3012), .Y(n2366) );
  MUX2X1 U7705 ( .B(arr[360]), .A(arr[401]), .S(n3012), .Y(n2365) );
  MUX2X1 U7706 ( .B(n2364), .A(n2361), .S(n3150), .Y(n2375) );
  MUX2X1 U7707 ( .B(arr[278]), .A(arr[319]), .S(n3012), .Y(n2369) );
  MUX2X1 U7708 ( .B(arr[196]), .A(arr[237]), .S(n3012), .Y(n2368) );
  MUX2X1 U7709 ( .B(arr[114]), .A(arr[155]), .S(n3012), .Y(n2372) );
  MUX2X1 U7710 ( .B(arr[32]), .A(arr[73]), .S(n3012), .Y(n2371) );
  MUX2X1 U7711 ( .B(n2370), .A(n2367), .S(n3150), .Y(n2374) );
  MUX2X1 U7712 ( .B(n2373), .A(n2358), .S(n3185), .Y(n2376) );
  MUX2X1 U7713 ( .B(arr[2575]), .A(arr[2616]), .S(n3012), .Y(n2380) );
  MUX2X1 U7714 ( .B(arr[2493]), .A(arr[2534]), .S(n3012), .Y(n2379) );
  MUX2X1 U7715 ( .B(arr[2411]), .A(arr[2452]), .S(n3012), .Y(n2383) );
  MUX2X1 U7716 ( .B(arr[2329]), .A(arr[2370]), .S(n3012), .Y(n2382) );
  MUX2X1 U7717 ( .B(n2381), .A(n2378), .S(n3150), .Y(n2392) );
  MUX2X1 U7718 ( .B(arr[2247]), .A(arr[2288]), .S(n3013), .Y(n2386) );
  MUX2X1 U7719 ( .B(arr[2165]), .A(arr[2206]), .S(n3013), .Y(n2385) );
  MUX2X1 U7720 ( .B(arr[2083]), .A(arr[2124]), .S(n3013), .Y(n2389) );
  MUX2X1 U7721 ( .B(arr[2001]), .A(arr[2042]), .S(n3013), .Y(n2388) );
  MUX2X1 U7722 ( .B(n2387), .A(n2384), .S(n3150), .Y(n2391) );
  MUX2X1 U7723 ( .B(arr[1919]), .A(arr[1960]), .S(n3013), .Y(n2395) );
  MUX2X1 U7724 ( .B(arr[1837]), .A(arr[1878]), .S(n3013), .Y(n2394) );
  MUX2X1 U7725 ( .B(arr[1755]), .A(arr[1796]), .S(n3013), .Y(n2398) );
  MUX2X1 U7726 ( .B(arr[1673]), .A(arr[1714]), .S(n3013), .Y(n2397) );
  MUX2X1 U7727 ( .B(n2396), .A(n2393), .S(n3150), .Y(n2407) );
  MUX2X1 U7728 ( .B(arr[1591]), .A(arr[1632]), .S(n3013), .Y(n2401) );
  MUX2X1 U7729 ( .B(arr[1509]), .A(arr[1550]), .S(n3013), .Y(n2400) );
  MUX2X1 U7730 ( .B(arr[1427]), .A(arr[1468]), .S(n3013), .Y(n2404) );
  MUX2X1 U7731 ( .B(arr[1345]), .A(arr[1386]), .S(n3013), .Y(n2403) );
  MUX2X1 U7732 ( .B(n2402), .A(n2399), .S(n3150), .Y(n2406) );
  MUX2X1 U7733 ( .B(n2405), .A(n2390), .S(n3185), .Y(n2439) );
  MUX2X1 U7734 ( .B(arr[1263]), .A(arr[1304]), .S(n3014), .Y(n2410) );
  MUX2X1 U7735 ( .B(arr[1181]), .A(arr[1222]), .S(n3014), .Y(n2409) );
  MUX2X1 U7736 ( .B(arr[1099]), .A(arr[1140]), .S(n3014), .Y(n2413) );
  MUX2X1 U7737 ( .B(arr[1017]), .A(arr[1058]), .S(n3014), .Y(n2412) );
  MUX2X1 U7738 ( .B(n2411), .A(n2408), .S(n3151), .Y(n2422) );
  MUX2X1 U7739 ( .B(arr[935]), .A(arr[976]), .S(n3014), .Y(n2416) );
  MUX2X1 U7740 ( .B(arr[853]), .A(arr[894]), .S(n3014), .Y(n2415) );
  MUX2X1 U7741 ( .B(arr[771]), .A(arr[812]), .S(n3014), .Y(n2419) );
  MUX2X1 U7742 ( .B(arr[689]), .A(arr[730]), .S(n3014), .Y(n2418) );
  MUX2X1 U7743 ( .B(n2417), .A(n2414), .S(n3151), .Y(n2421) );
  MUX2X1 U7744 ( .B(arr[607]), .A(arr[648]), .S(n3014), .Y(n2425) );
  MUX2X1 U7745 ( .B(arr[525]), .A(arr[566]), .S(n3014), .Y(n2424) );
  MUX2X1 U7746 ( .B(arr[443]), .A(arr[484]), .S(n3014), .Y(n2428) );
  MUX2X1 U7747 ( .B(arr[361]), .A(arr[402]), .S(n3014), .Y(n2427) );
  MUX2X1 U7748 ( .B(n2426), .A(n2423), .S(n3151), .Y(n2437) );
  MUX2X1 U7749 ( .B(arr[279]), .A(arr[320]), .S(n3015), .Y(n2431) );
  MUX2X1 U7750 ( .B(arr[197]), .A(arr[238]), .S(n3015), .Y(n2430) );
  MUX2X1 U7751 ( .B(arr[115]), .A(arr[156]), .S(n3015), .Y(n2434) );
  MUX2X1 U7752 ( .B(arr[33]), .A(arr[74]), .S(n3015), .Y(n2433) );
  MUX2X1 U7753 ( .B(n2432), .A(n2429), .S(n3151), .Y(n2436) );
  MUX2X1 U7754 ( .B(n2435), .A(n2420), .S(n3185), .Y(n2438) );
  MUX2X1 U7755 ( .B(arr[2576]), .A(arr[2617]), .S(n3015), .Y(n2442) );
  MUX2X1 U7756 ( .B(arr[2494]), .A(arr[2535]), .S(n3015), .Y(n2441) );
  MUX2X1 U7757 ( .B(arr[2412]), .A(arr[2453]), .S(n3015), .Y(n2445) );
  MUX2X1 U7758 ( .B(arr[2330]), .A(arr[2371]), .S(n3015), .Y(n2444) );
  MUX2X1 U7759 ( .B(n2443), .A(n2440), .S(n3151), .Y(n2454) );
  MUX2X1 U7760 ( .B(arr[2248]), .A(arr[2289]), .S(n3015), .Y(n2448) );
  MUX2X1 U7761 ( .B(arr[2166]), .A(arr[2207]), .S(n3015), .Y(n2447) );
  MUX2X1 U7762 ( .B(arr[2084]), .A(arr[2125]), .S(n3015), .Y(n2451) );
  MUX2X1 U7763 ( .B(arr[2002]), .A(arr[2043]), .S(n3015), .Y(n2450) );
  MUX2X1 U7764 ( .B(n2449), .A(n2446), .S(n3151), .Y(n2453) );
  MUX2X1 U7765 ( .B(arr[1920]), .A(arr[1961]), .S(n3016), .Y(n2457) );
  MUX2X1 U7766 ( .B(arr[1838]), .A(arr[1879]), .S(n3016), .Y(n2456) );
  MUX2X1 U7767 ( .B(arr[1756]), .A(arr[1797]), .S(n3016), .Y(n2460) );
  MUX2X1 U7768 ( .B(arr[1674]), .A(arr[1715]), .S(n3016), .Y(n2459) );
  MUX2X1 U7769 ( .B(n2458), .A(n2455), .S(n3151), .Y(n2469) );
  MUX2X1 U7770 ( .B(arr[1592]), .A(arr[1633]), .S(n3016), .Y(n2463) );
  MUX2X1 U7771 ( .B(arr[1510]), .A(arr[1551]), .S(n3016), .Y(n2462) );
  MUX2X1 U7772 ( .B(arr[1428]), .A(arr[1469]), .S(n3016), .Y(n2466) );
  MUX2X1 U7773 ( .B(arr[1346]), .A(arr[1387]), .S(n3016), .Y(n2465) );
  MUX2X1 U7774 ( .B(n2464), .A(n2461), .S(n3151), .Y(n2468) );
  MUX2X1 U7775 ( .B(n2467), .A(n2452), .S(n3185), .Y(n2501) );
  MUX2X1 U7776 ( .B(arr[1264]), .A(arr[1305]), .S(n3016), .Y(n2472) );
  MUX2X1 U7777 ( .B(arr[1182]), .A(arr[1223]), .S(n3016), .Y(n2471) );
  MUX2X1 U7778 ( .B(arr[1100]), .A(arr[1141]), .S(n3016), .Y(n2475) );
  MUX2X1 U7779 ( .B(arr[1018]), .A(arr[1059]), .S(n3016), .Y(n2474) );
  MUX2X1 U7780 ( .B(n2473), .A(n2470), .S(n3151), .Y(n2484) );
  MUX2X1 U7781 ( .B(arr[936]), .A(arr[977]), .S(n3017), .Y(n2478) );
  MUX2X1 U7782 ( .B(arr[854]), .A(arr[895]), .S(n3017), .Y(n2477) );
  MUX2X1 U7783 ( .B(arr[772]), .A(arr[813]), .S(n3017), .Y(n2481) );
  MUX2X1 U7784 ( .B(arr[690]), .A(arr[731]), .S(n3017), .Y(n2480) );
  MUX2X1 U7785 ( .B(n2479), .A(n2476), .S(n3151), .Y(n2483) );
  MUX2X1 U7786 ( .B(arr[608]), .A(arr[649]), .S(n3017), .Y(n2487) );
  MUX2X1 U7787 ( .B(arr[526]), .A(arr[567]), .S(n3017), .Y(n2486) );
  MUX2X1 U7788 ( .B(arr[444]), .A(arr[485]), .S(n3017), .Y(n2490) );
  MUX2X1 U7789 ( .B(arr[362]), .A(arr[403]), .S(n3017), .Y(n2489) );
  MUX2X1 U7790 ( .B(n2488), .A(n2485), .S(n3151), .Y(n2499) );
  MUX2X1 U7791 ( .B(arr[280]), .A(arr[321]), .S(n3017), .Y(n2493) );
  MUX2X1 U7792 ( .B(arr[198]), .A(arr[239]), .S(n3017), .Y(n2492) );
  MUX2X1 U7793 ( .B(arr[116]), .A(arr[157]), .S(n3017), .Y(n2496) );
  MUX2X1 U7794 ( .B(arr[34]), .A(arr[75]), .S(n3017), .Y(n2495) );
  MUX2X1 U7795 ( .B(n2494), .A(n2491), .S(n3151), .Y(n2498) );
  MUX2X1 U7796 ( .B(n2497), .A(n2482), .S(n3185), .Y(n2500) );
  MUX2X1 U7797 ( .B(arr[2577]), .A(arr[2618]), .S(n3018), .Y(n2504) );
  MUX2X1 U7798 ( .B(arr[2495]), .A(arr[2536]), .S(n3018), .Y(n2503) );
  MUX2X1 U7799 ( .B(arr[2413]), .A(arr[2454]), .S(n3018), .Y(n2507) );
  MUX2X1 U7800 ( .B(arr[2331]), .A(arr[2372]), .S(n3018), .Y(n2506) );
  MUX2X1 U7801 ( .B(n2505), .A(n2502), .S(n3152), .Y(n2516) );
  MUX2X1 U7802 ( .B(arr[2249]), .A(arr[2290]), .S(n3018), .Y(n2510) );
  MUX2X1 U7803 ( .B(arr[2167]), .A(arr[2208]), .S(n3018), .Y(n2509) );
  MUX2X1 U7804 ( .B(arr[2085]), .A(arr[2126]), .S(n3018), .Y(n2513) );
  MUX2X1 U7805 ( .B(arr[2003]), .A(arr[2044]), .S(n3018), .Y(n2512) );
  MUX2X1 U7806 ( .B(n2511), .A(n2508), .S(n3152), .Y(n2515) );
  MUX2X1 U7807 ( .B(arr[1921]), .A(arr[1962]), .S(n3018), .Y(n2519) );
  MUX2X1 U7808 ( .B(arr[1839]), .A(arr[1880]), .S(n3018), .Y(n2518) );
  MUX2X1 U7809 ( .B(arr[1757]), .A(arr[1798]), .S(n3018), .Y(n2522) );
  MUX2X1 U7810 ( .B(arr[1675]), .A(arr[1716]), .S(n3018), .Y(n2521) );
  MUX2X1 U7811 ( .B(n2520), .A(n2517), .S(n3152), .Y(n2531) );
  MUX2X1 U7812 ( .B(arr[1593]), .A(arr[1634]), .S(n3019), .Y(n2525) );
  MUX2X1 U7813 ( .B(arr[1511]), .A(arr[1552]), .S(n3019), .Y(n2524) );
  MUX2X1 U7814 ( .B(arr[1429]), .A(arr[1470]), .S(n3019), .Y(n2528) );
  MUX2X1 U7815 ( .B(arr[1347]), .A(arr[1388]), .S(n3019), .Y(n2527) );
  MUX2X1 U7816 ( .B(n2526), .A(n2523), .S(n3152), .Y(n2530) );
  MUX2X1 U7817 ( .B(n2529), .A(n2514), .S(n3186), .Y(n2563) );
  MUX2X1 U7818 ( .B(arr[1265]), .A(arr[1306]), .S(n3019), .Y(n2534) );
  MUX2X1 U7819 ( .B(arr[1183]), .A(arr[1224]), .S(n3019), .Y(n2533) );
  MUX2X1 U7820 ( .B(arr[1101]), .A(arr[1142]), .S(n3019), .Y(n2537) );
  MUX2X1 U7821 ( .B(arr[1019]), .A(arr[1060]), .S(n3019), .Y(n2536) );
  MUX2X1 U7822 ( .B(n2535), .A(n2532), .S(n3152), .Y(n2546) );
  MUX2X1 U7823 ( .B(arr[937]), .A(arr[978]), .S(n3019), .Y(n2540) );
  MUX2X1 U7824 ( .B(arr[855]), .A(arr[896]), .S(n3019), .Y(n2539) );
  MUX2X1 U7825 ( .B(arr[773]), .A(arr[814]), .S(n3019), .Y(n2543) );
  MUX2X1 U7826 ( .B(arr[691]), .A(arr[732]), .S(n3019), .Y(n2542) );
  MUX2X1 U7827 ( .B(n2541), .A(n2538), .S(n3152), .Y(n2545) );
  MUX2X1 U7828 ( .B(arr[609]), .A(arr[650]), .S(n3020), .Y(n2549) );
  MUX2X1 U7829 ( .B(arr[527]), .A(arr[568]), .S(n3020), .Y(n2548) );
  MUX2X1 U7830 ( .B(arr[445]), .A(arr[486]), .S(n3020), .Y(n2552) );
  MUX2X1 U7831 ( .B(arr[363]), .A(arr[404]), .S(n3020), .Y(n2551) );
  MUX2X1 U7832 ( .B(n2550), .A(n2547), .S(n3152), .Y(n2561) );
  MUX2X1 U7833 ( .B(arr[281]), .A(arr[322]), .S(n3020), .Y(n2555) );
  MUX2X1 U7834 ( .B(arr[199]), .A(arr[240]), .S(n3020), .Y(n2554) );
  MUX2X1 U7835 ( .B(arr[117]), .A(arr[158]), .S(n3020), .Y(n2558) );
  MUX2X1 U7836 ( .B(arr[35]), .A(arr[76]), .S(n3020), .Y(n2557) );
  MUX2X1 U7837 ( .B(n2556), .A(n2553), .S(n3152), .Y(n2560) );
  MUX2X1 U7838 ( .B(n2559), .A(n2544), .S(n3186), .Y(n2562) );
  MUX2X1 U7839 ( .B(arr[2578]), .A(arr[2619]), .S(n3020), .Y(n2566) );
  MUX2X1 U7840 ( .B(arr[2496]), .A(arr[2537]), .S(n3020), .Y(n2565) );
  MUX2X1 U7841 ( .B(arr[2414]), .A(arr[2455]), .S(n3020), .Y(n2569) );
  MUX2X1 U7842 ( .B(arr[2332]), .A(arr[2373]), .S(n3020), .Y(n2568) );
  MUX2X1 U7843 ( .B(n2567), .A(n2564), .S(n3152), .Y(n2578) );
  MUX2X1 U7844 ( .B(arr[2250]), .A(arr[2291]), .S(n3021), .Y(n2572) );
  MUX2X1 U7845 ( .B(arr[2168]), .A(arr[2209]), .S(n3021), .Y(n2571) );
  MUX2X1 U7846 ( .B(arr[2086]), .A(arr[2127]), .S(n3021), .Y(n2575) );
  MUX2X1 U7847 ( .B(arr[2004]), .A(arr[2045]), .S(n3021), .Y(n2574) );
  MUX2X1 U7848 ( .B(n2573), .A(n2570), .S(n3152), .Y(n2577) );
  MUX2X1 U7849 ( .B(arr[1922]), .A(arr[1963]), .S(n3021), .Y(n2581) );
  MUX2X1 U7850 ( .B(arr[1840]), .A(arr[1881]), .S(n3021), .Y(n2580) );
  MUX2X1 U7851 ( .B(arr[1758]), .A(arr[1799]), .S(n3021), .Y(n2584) );
  MUX2X1 U7852 ( .B(arr[1676]), .A(arr[1717]), .S(n3021), .Y(n2583) );
  MUX2X1 U7853 ( .B(n2582), .A(n2579), .S(n3152), .Y(n2593) );
  MUX2X1 U7854 ( .B(arr[1594]), .A(arr[1635]), .S(n3021), .Y(n2587) );
  MUX2X1 U7855 ( .B(arr[1512]), .A(arr[1553]), .S(n3021), .Y(n2586) );
  MUX2X1 U7856 ( .B(arr[1430]), .A(arr[1471]), .S(n3021), .Y(n2590) );
  MUX2X1 U7857 ( .B(arr[1348]), .A(arr[1389]), .S(n3021), .Y(n2589) );
  MUX2X1 U7858 ( .B(n2588), .A(n2585), .S(n3152), .Y(n2592) );
  MUX2X1 U7859 ( .B(n2591), .A(n2576), .S(n3186), .Y(n2625) );
  MUX2X1 U7860 ( .B(arr[1266]), .A(arr[1307]), .S(n3022), .Y(n2596) );
  MUX2X1 U7861 ( .B(arr[1184]), .A(arr[1225]), .S(n3022), .Y(n2595) );
  MUX2X1 U7862 ( .B(arr[1102]), .A(arr[1143]), .S(n3022), .Y(n2599) );
  MUX2X1 U7863 ( .B(arr[1020]), .A(arr[1061]), .S(n3022), .Y(n2598) );
  MUX2X1 U7864 ( .B(n2597), .A(n2594), .S(n3153), .Y(n2608) );
  MUX2X1 U7865 ( .B(arr[938]), .A(arr[979]), .S(n3022), .Y(n2602) );
  MUX2X1 U7866 ( .B(arr[856]), .A(arr[897]), .S(n3022), .Y(n2601) );
  MUX2X1 U7867 ( .B(arr[774]), .A(arr[815]), .S(n3022), .Y(n2605) );
  MUX2X1 U7868 ( .B(arr[692]), .A(arr[733]), .S(n3022), .Y(n2604) );
  MUX2X1 U7869 ( .B(n2603), .A(n2600), .S(n3153), .Y(n2607) );
  MUX2X1 U7870 ( .B(arr[610]), .A(arr[651]), .S(n3022), .Y(n2611) );
  MUX2X1 U7871 ( .B(arr[528]), .A(arr[569]), .S(n3022), .Y(n2610) );
  MUX2X1 U7872 ( .B(arr[446]), .A(arr[487]), .S(n3022), .Y(n2614) );
  MUX2X1 U7873 ( .B(arr[364]), .A(arr[405]), .S(n3022), .Y(n2613) );
  MUX2X1 U7874 ( .B(n2612), .A(n2609), .S(n3153), .Y(n2623) );
  MUX2X1 U7875 ( .B(arr[282]), .A(arr[323]), .S(n3023), .Y(n2617) );
  MUX2X1 U7876 ( .B(arr[200]), .A(arr[241]), .S(n3023), .Y(n2616) );
  MUX2X1 U7877 ( .B(arr[118]), .A(arr[159]), .S(n3023), .Y(n2620) );
  MUX2X1 U7878 ( .B(arr[36]), .A(arr[77]), .S(n3023), .Y(n2619) );
  MUX2X1 U7879 ( .B(n2618), .A(n2615), .S(n3153), .Y(n2622) );
  MUX2X1 U7880 ( .B(n2621), .A(n2606), .S(n3186), .Y(n2624) );
  MUX2X1 U7881 ( .B(arr[2579]), .A(arr[2620]), .S(n3023), .Y(n2628) );
  MUX2X1 U7882 ( .B(arr[2497]), .A(arr[2538]), .S(n3023), .Y(n2627) );
  MUX2X1 U7883 ( .B(arr[2415]), .A(arr[2456]), .S(n3023), .Y(n2631) );
  MUX2X1 U7884 ( .B(arr[2333]), .A(arr[2374]), .S(n3023), .Y(n2630) );
  MUX2X1 U7885 ( .B(n2629), .A(n2626), .S(n3153), .Y(n2640) );
  MUX2X1 U7886 ( .B(arr[2251]), .A(arr[2292]), .S(n3023), .Y(n2634) );
  MUX2X1 U7887 ( .B(arr[2169]), .A(arr[2210]), .S(n3023), .Y(n2633) );
  MUX2X1 U7888 ( .B(arr[2087]), .A(arr[2128]), .S(n3023), .Y(n2637) );
  MUX2X1 U7889 ( .B(arr[2005]), .A(arr[2046]), .S(n3023), .Y(n2636) );
  MUX2X1 U7890 ( .B(n2635), .A(n2632), .S(n3153), .Y(n2639) );
  MUX2X1 U7891 ( .B(arr[1923]), .A(arr[1964]), .S(n3024), .Y(n2643) );
  MUX2X1 U7892 ( .B(arr[1841]), .A(arr[1882]), .S(n3024), .Y(n2642) );
  MUX2X1 U7893 ( .B(arr[1759]), .A(arr[1800]), .S(n3024), .Y(n2646) );
  MUX2X1 U7894 ( .B(arr[1677]), .A(arr[1718]), .S(n3024), .Y(n2645) );
  MUX2X1 U7895 ( .B(n2644), .A(n2641), .S(n3153), .Y(n2655) );
  MUX2X1 U7896 ( .B(arr[1595]), .A(arr[1636]), .S(n3024), .Y(n2649) );
  MUX2X1 U7897 ( .B(arr[1513]), .A(arr[1554]), .S(n3024), .Y(n2648) );
  MUX2X1 U7898 ( .B(arr[1431]), .A(arr[1472]), .S(n3024), .Y(n2652) );
  MUX2X1 U7899 ( .B(arr[1349]), .A(arr[1390]), .S(n3024), .Y(n2651) );
  MUX2X1 U7900 ( .B(n2650), .A(n2647), .S(n3153), .Y(n2654) );
  MUX2X1 U7901 ( .B(n2653), .A(n2638), .S(n3186), .Y(n2687) );
  MUX2X1 U7902 ( .B(arr[1267]), .A(arr[1308]), .S(n3024), .Y(n2658) );
  MUX2X1 U7903 ( .B(arr[1185]), .A(arr[1226]), .S(n3024), .Y(n2657) );
  MUX2X1 U7904 ( .B(arr[1103]), .A(arr[1144]), .S(n3024), .Y(n2661) );
  MUX2X1 U7905 ( .B(arr[1021]), .A(arr[1062]), .S(n3024), .Y(n2660) );
  MUX2X1 U7906 ( .B(n2659), .A(n2656), .S(n3153), .Y(n2670) );
  MUX2X1 U7907 ( .B(arr[939]), .A(arr[980]), .S(n3025), .Y(n2664) );
  MUX2X1 U7908 ( .B(arr[857]), .A(arr[898]), .S(n3025), .Y(n2663) );
  MUX2X1 U7909 ( .B(arr[775]), .A(arr[816]), .S(n3025), .Y(n2667) );
  MUX2X1 U7910 ( .B(arr[693]), .A(arr[734]), .S(n3025), .Y(n2666) );
  MUX2X1 U7911 ( .B(n2665), .A(n2662), .S(n3153), .Y(n2669) );
  MUX2X1 U7912 ( .B(arr[611]), .A(arr[652]), .S(n3025), .Y(n2673) );
  MUX2X1 U7913 ( .B(arr[529]), .A(arr[570]), .S(n3025), .Y(n2672) );
  MUX2X1 U7914 ( .B(arr[447]), .A(arr[488]), .S(n3025), .Y(n2676) );
  MUX2X1 U7915 ( .B(arr[365]), .A(arr[406]), .S(n3025), .Y(n2675) );
  MUX2X1 U7916 ( .B(n2674), .A(n2671), .S(n3153), .Y(n2685) );
  MUX2X1 U7917 ( .B(arr[283]), .A(arr[324]), .S(n3025), .Y(n2679) );
  MUX2X1 U7918 ( .B(arr[201]), .A(arr[242]), .S(n3025), .Y(n2678) );
  MUX2X1 U7919 ( .B(arr[119]), .A(arr[160]), .S(n3025), .Y(n2682) );
  MUX2X1 U7920 ( .B(arr[37]), .A(arr[78]), .S(n3025), .Y(n2681) );
  MUX2X1 U7921 ( .B(n2680), .A(n2677), .S(n3153), .Y(n2684) );
  MUX2X1 U7922 ( .B(n2683), .A(n2668), .S(n3186), .Y(n2686) );
  MUX2X1 U7923 ( .B(arr[2580]), .A(arr[2621]), .S(n3026), .Y(n2690) );
  MUX2X1 U7924 ( .B(arr[2498]), .A(arr[2539]), .S(n3026), .Y(n2689) );
  MUX2X1 U7925 ( .B(arr[2416]), .A(arr[2457]), .S(n3026), .Y(n2693) );
  MUX2X1 U7926 ( .B(arr[2334]), .A(arr[2375]), .S(n3026), .Y(n2692) );
  MUX2X1 U7927 ( .B(n2691), .A(n2688), .S(n3154), .Y(n2702) );
  MUX2X1 U7928 ( .B(arr[2252]), .A(arr[2293]), .S(n3026), .Y(n2696) );
  MUX2X1 U7929 ( .B(arr[2170]), .A(arr[2211]), .S(n3026), .Y(n2695) );
  MUX2X1 U7930 ( .B(arr[2088]), .A(arr[2129]), .S(n3026), .Y(n2699) );
  MUX2X1 U7931 ( .B(arr[2006]), .A(arr[2047]), .S(n3026), .Y(n2698) );
  MUX2X1 U7932 ( .B(n2697), .A(n2694), .S(n3154), .Y(n2701) );
  MUX2X1 U7933 ( .B(arr[1924]), .A(arr[1965]), .S(n3026), .Y(n2705) );
  MUX2X1 U7934 ( .B(arr[1842]), .A(arr[1883]), .S(n3026), .Y(n2704) );
  MUX2X1 U7935 ( .B(arr[1760]), .A(arr[1801]), .S(n3026), .Y(n2708) );
  MUX2X1 U7936 ( .B(arr[1678]), .A(arr[1719]), .S(n3026), .Y(n2707) );
  MUX2X1 U7937 ( .B(n2706), .A(n2703), .S(n3154), .Y(n2717) );
  MUX2X1 U7938 ( .B(arr[1596]), .A(arr[1637]), .S(n3027), .Y(n2711) );
  MUX2X1 U7939 ( .B(arr[1514]), .A(arr[1555]), .S(n3027), .Y(n2710) );
  MUX2X1 U7940 ( .B(arr[1432]), .A(arr[1473]), .S(n3027), .Y(n2714) );
  MUX2X1 U7941 ( .B(arr[1350]), .A(arr[1391]), .S(n3027), .Y(n2713) );
  MUX2X1 U7942 ( .B(n2712), .A(n2709), .S(n3154), .Y(n2716) );
  MUX2X1 U7943 ( .B(n2715), .A(n2700), .S(n3186), .Y(n2762) );
  MUX2X1 U7944 ( .B(arr[1268]), .A(arr[1309]), .S(n3027), .Y(n2720) );
  MUX2X1 U7945 ( .B(arr[1186]), .A(arr[1227]), .S(n3027), .Y(n2719) );
  MUX2X1 U7946 ( .B(arr[1104]), .A(arr[1145]), .S(n3027), .Y(n2723) );
  MUX2X1 U7947 ( .B(arr[1022]), .A(arr[1063]), .S(n3027), .Y(n2722) );
  MUX2X1 U7948 ( .B(n2721), .A(n2718), .S(n3154), .Y(n2745) );
  MUX2X1 U7949 ( .B(arr[940]), .A(arr[981]), .S(n3027), .Y(n2739) );
  MUX2X1 U7950 ( .B(arr[858]), .A(arr[899]), .S(n3027), .Y(n2738) );
  MUX2X1 U7951 ( .B(arr[776]), .A(arr[817]), .S(n3027), .Y(n2742) );
  MUX2X1 U7952 ( .B(arr[694]), .A(arr[735]), .S(n3027), .Y(n2741) );
  MUX2X1 U7953 ( .B(n2740), .A(n2724), .S(n3154), .Y(n2744) );
  MUX2X1 U7954 ( .B(arr[612]), .A(arr[653]), .S(n3028), .Y(n2748) );
  MUX2X1 U7955 ( .B(arr[530]), .A(arr[571]), .S(n3028), .Y(n2747) );
  MUX2X1 U7956 ( .B(arr[448]), .A(arr[489]), .S(n3028), .Y(n2751) );
  MUX2X1 U7957 ( .B(arr[366]), .A(arr[407]), .S(n3028), .Y(n2750) );
  MUX2X1 U7958 ( .B(n2749), .A(n2746), .S(n3154), .Y(n2760) );
  MUX2X1 U7959 ( .B(arr[284]), .A(arr[325]), .S(n3028), .Y(n2754) );
  MUX2X1 U7960 ( .B(arr[202]), .A(arr[243]), .S(n3028), .Y(n2753) );
  MUX2X1 U7961 ( .B(arr[120]), .A(arr[161]), .S(n3028), .Y(n2757) );
  MUX2X1 U7962 ( .B(arr[38]), .A(arr[79]), .S(n3028), .Y(n2756) );
  MUX2X1 U7963 ( .B(n2755), .A(n2752), .S(n3154), .Y(n2759) );
  MUX2X1 U7964 ( .B(n2758), .A(n2743), .S(n3186), .Y(n2761) );
  MUX2X1 U7965 ( .B(arr[2581]), .A(arr[2622]), .S(n3028), .Y(n2765) );
  MUX2X1 U7966 ( .B(arr[2499]), .A(arr[2540]), .S(n3028), .Y(n2764) );
  MUX2X1 U7967 ( .B(arr[2417]), .A(arr[2458]), .S(n3028), .Y(n2768) );
  MUX2X1 U7968 ( .B(arr[2335]), .A(arr[2376]), .S(n3028), .Y(n2767) );
  MUX2X1 U7969 ( .B(n2766), .A(n2763), .S(n3154), .Y(n2777) );
  MUX2X1 U7970 ( .B(arr[2253]), .A(arr[2294]), .S(n3029), .Y(n2771) );
  MUX2X1 U7971 ( .B(arr[2171]), .A(arr[2212]), .S(n3029), .Y(n2770) );
  MUX2X1 U7972 ( .B(arr[2089]), .A(arr[2130]), .S(n3029), .Y(n2774) );
  MUX2X1 U7973 ( .B(arr[2007]), .A(arr[2048]), .S(n3029), .Y(n2773) );
  MUX2X1 U7974 ( .B(n2772), .A(n2769), .S(n3154), .Y(n2776) );
  MUX2X1 U7975 ( .B(arr[1925]), .A(arr[1966]), .S(n3029), .Y(n2780) );
  MUX2X1 U7976 ( .B(arr[1843]), .A(arr[1884]), .S(n3029), .Y(n2779) );
  MUX2X1 U7977 ( .B(arr[1761]), .A(arr[1802]), .S(n3029), .Y(n2783) );
  MUX2X1 U7978 ( .B(arr[1679]), .A(arr[1720]), .S(n3029), .Y(n2782) );
  MUX2X1 U7979 ( .B(n2781), .A(n2778), .S(n3154), .Y(n2792) );
  MUX2X1 U7980 ( .B(arr[1597]), .A(arr[1638]), .S(n3029), .Y(n2786) );
  MUX2X1 U7981 ( .B(arr[1515]), .A(arr[1556]), .S(n3029), .Y(n2785) );
  MUX2X1 U7982 ( .B(arr[1433]), .A(arr[1474]), .S(n3029), .Y(n2789) );
  MUX2X1 U7983 ( .B(arr[1351]), .A(arr[1392]), .S(n3029), .Y(n2788) );
  MUX2X1 U7984 ( .B(n2787), .A(n2784), .S(n3154), .Y(n2791) );
  MUX2X1 U7985 ( .B(n2790), .A(n2775), .S(n3186), .Y(n2824) );
  MUX2X1 U7986 ( .B(arr[1269]), .A(arr[1310]), .S(n3030), .Y(n2795) );
  MUX2X1 U7987 ( .B(arr[1187]), .A(arr[1228]), .S(n3030), .Y(n2794) );
  MUX2X1 U7988 ( .B(arr[1105]), .A(arr[1146]), .S(n3030), .Y(n2798) );
  MUX2X1 U7989 ( .B(arr[1023]), .A(arr[1064]), .S(n3030), .Y(n2797) );
  MUX2X1 U7990 ( .B(n2796), .A(n2793), .S(n3155), .Y(n2807) );
  MUX2X1 U7991 ( .B(arr[941]), .A(arr[982]), .S(n3030), .Y(n2801) );
  MUX2X1 U7992 ( .B(arr[859]), .A(arr[900]), .S(n3030), .Y(n2800) );
  MUX2X1 U7993 ( .B(arr[777]), .A(arr[818]), .S(n3030), .Y(n2804) );
  MUX2X1 U7994 ( .B(arr[695]), .A(arr[736]), .S(n3030), .Y(n2803) );
  MUX2X1 U7995 ( .B(n2802), .A(n2799), .S(n3155), .Y(n2806) );
  MUX2X1 U7996 ( .B(arr[613]), .A(arr[654]), .S(n3030), .Y(n2810) );
  MUX2X1 U7997 ( .B(arr[531]), .A(arr[572]), .S(n3030), .Y(n2809) );
  MUX2X1 U7998 ( .B(arr[449]), .A(arr[490]), .S(n3030), .Y(n2813) );
  MUX2X1 U7999 ( .B(arr[367]), .A(arr[408]), .S(n3030), .Y(n2812) );
  MUX2X1 U8000 ( .B(n2811), .A(n2808), .S(n3155), .Y(n2822) );
  MUX2X1 U8001 ( .B(arr[285]), .A(arr[326]), .S(n3031), .Y(n2816) );
  MUX2X1 U8002 ( .B(arr[203]), .A(arr[244]), .S(n3031), .Y(n2815) );
  MUX2X1 U8003 ( .B(arr[121]), .A(arr[162]), .S(n3031), .Y(n2819) );
  MUX2X1 U8004 ( .B(arr[39]), .A(arr[80]), .S(n3031), .Y(n2818) );
  MUX2X1 U8005 ( .B(n2817), .A(n2814), .S(n3155), .Y(n2821) );
  MUX2X1 U8006 ( .B(n2820), .A(n2805), .S(n3186), .Y(n2823) );
  MUX2X1 U8007 ( .B(arr[2582]), .A(arr[2623]), .S(n3031), .Y(n2827) );
  MUX2X1 U8008 ( .B(arr[2500]), .A(arr[2541]), .S(n3031), .Y(n2826) );
  MUX2X1 U8009 ( .B(arr[2418]), .A(arr[2459]), .S(n3031), .Y(n2830) );
  MUX2X1 U8010 ( .B(arr[2336]), .A(arr[2377]), .S(n3031), .Y(n2829) );
  MUX2X1 U8011 ( .B(n2828), .A(n2825), .S(n3155), .Y(n2839) );
  MUX2X1 U8012 ( .B(arr[2254]), .A(arr[2295]), .S(n3031), .Y(n2833) );
  MUX2X1 U8013 ( .B(arr[2172]), .A(arr[2213]), .S(n3031), .Y(n2832) );
  MUX2X1 U8014 ( .B(arr[2090]), .A(arr[2131]), .S(n3031), .Y(n2836) );
  MUX2X1 U8015 ( .B(arr[2008]), .A(arr[2049]), .S(n3031), .Y(n2835) );
  MUX2X1 U8016 ( .B(n2834), .A(n2831), .S(n3155), .Y(n2838) );
  MUX2X1 U8017 ( .B(arr[1926]), .A(arr[1967]), .S(n3032), .Y(n2842) );
  MUX2X1 U8018 ( .B(arr[1844]), .A(arr[1885]), .S(n3032), .Y(n2841) );
  MUX2X1 U8019 ( .B(arr[1762]), .A(arr[1803]), .S(n3032), .Y(n2845) );
  MUX2X1 U8020 ( .B(arr[1680]), .A(arr[1721]), .S(n3032), .Y(n2844) );
  MUX2X1 U8021 ( .B(n2843), .A(n2840), .S(n3155), .Y(n2854) );
  MUX2X1 U8022 ( .B(arr[1598]), .A(arr[1639]), .S(n3032), .Y(n2848) );
  MUX2X1 U8023 ( .B(arr[1516]), .A(arr[1557]), .S(n3032), .Y(n2847) );
  MUX2X1 U8024 ( .B(arr[1434]), .A(arr[1475]), .S(n3032), .Y(n2851) );
  MUX2X1 U8025 ( .B(arr[1352]), .A(arr[1393]), .S(n3032), .Y(n2850) );
  MUX2X1 U8026 ( .B(n2849), .A(n2846), .S(n3155), .Y(n2853) );
  MUX2X1 U8027 ( .B(n2852), .A(n2837), .S(n3186), .Y(n2886) );
  MUX2X1 U8028 ( .B(arr[1270]), .A(arr[1311]), .S(n3032), .Y(n2857) );
  MUX2X1 U8029 ( .B(arr[1188]), .A(arr[1229]), .S(n3032), .Y(n2856) );
  MUX2X1 U8030 ( .B(arr[1106]), .A(arr[1147]), .S(n3032), .Y(n2860) );
  MUX2X1 U8031 ( .B(arr[1024]), .A(arr[1065]), .S(n3032), .Y(n2859) );
  MUX2X1 U8032 ( .B(n2858), .A(n2855), .S(n3155), .Y(n2869) );
  MUX2X1 U8033 ( .B(arr[942]), .A(arr[983]), .S(n3033), .Y(n2863) );
  MUX2X1 U8034 ( .B(arr[860]), .A(arr[901]), .S(n3033), .Y(n2862) );
  MUX2X1 U8035 ( .B(arr[778]), .A(arr[819]), .S(n3033), .Y(n2866) );
  MUX2X1 U8036 ( .B(arr[696]), .A(arr[737]), .S(n3033), .Y(n2865) );
  MUX2X1 U8037 ( .B(n2864), .A(n2861), .S(n3155), .Y(n2868) );
  MUX2X1 U8038 ( .B(arr[614]), .A(arr[655]), .S(n3033), .Y(n2872) );
  MUX2X1 U8039 ( .B(arr[532]), .A(arr[573]), .S(n3033), .Y(n2871) );
  MUX2X1 U8040 ( .B(arr[450]), .A(arr[491]), .S(n3033), .Y(n2875) );
  MUX2X1 U8041 ( .B(arr[368]), .A(arr[409]), .S(n3033), .Y(n2874) );
  MUX2X1 U8042 ( .B(n2873), .A(n2870), .S(n3155), .Y(n2884) );
  MUX2X1 U8043 ( .B(arr[286]), .A(arr[327]), .S(n3033), .Y(n2878) );
  MUX2X1 U8044 ( .B(arr[204]), .A(arr[245]), .S(n3033), .Y(n2877) );
  MUX2X1 U8045 ( .B(arr[122]), .A(arr[163]), .S(n3033), .Y(n2881) );
  MUX2X1 U8046 ( .B(arr[40]), .A(arr[81]), .S(n3033), .Y(n2880) );
  MUX2X1 U8047 ( .B(n2879), .A(n2876), .S(n3155), .Y(n2883) );
  MUX2X1 U8048 ( .B(n2882), .A(n2867), .S(n3186), .Y(n2885) );
  BUFX2 U8049 ( .A(n6173), .Y(n3464) );
  BUFX2 U8050 ( .A(n6173), .Y(n3461) );
  BUFX2 U8051 ( .A(n6173), .Y(n3460) );
  BUFX2 U8052 ( .A(n6173), .Y(n3459) );
  BUFX2 U8053 ( .A(n6131), .Y(n3465) );
  BUFX2 U8054 ( .A(n6131), .Y(n3466) );
  BUFX2 U8055 ( .A(n6131), .Y(n3467) );
  BUFX2 U8056 ( .A(n6131), .Y(n3470) );
  BUFX2 U8057 ( .A(n6089), .Y(n3476) );
  BUFX2 U8058 ( .A(n6089), .Y(n3473) );
  BUFX2 U8059 ( .A(n6089), .Y(n3472) );
  BUFX2 U8060 ( .A(n6089), .Y(n3471) );
  BUFX2 U8061 ( .A(n6046), .Y(n3477) );
  BUFX2 U8062 ( .A(n6046), .Y(n3478) );
  BUFX2 U8063 ( .A(n6046), .Y(n3479) );
  BUFX2 U8064 ( .A(n6046), .Y(n3482) );
  BUFX2 U8065 ( .A(n6003), .Y(n3488) );
  BUFX2 U8066 ( .A(n6003), .Y(n3485) );
  BUFX2 U8067 ( .A(n6003), .Y(n3484) );
  BUFX2 U8068 ( .A(n6003), .Y(n3483) );
  BUFX2 U8069 ( .A(n5961), .Y(n3489) );
  BUFX2 U8070 ( .A(n5961), .Y(n3490) );
  BUFX2 U8071 ( .A(n5961), .Y(n3491) );
  BUFX2 U8072 ( .A(n5961), .Y(n3494) );
  BUFX2 U8073 ( .A(n5919), .Y(n3500) );
  BUFX2 U8074 ( .A(n5919), .Y(n3497) );
  BUFX2 U8075 ( .A(n5919), .Y(n3496) );
  BUFX2 U8076 ( .A(n5919), .Y(n3495) );
  BUFX2 U8077 ( .A(n5876), .Y(n3501) );
  BUFX2 U8078 ( .A(n5876), .Y(n3502) );
  BUFX2 U8079 ( .A(n5876), .Y(n3503) );
  BUFX2 U8080 ( .A(n5876), .Y(n3506) );
  BUFX2 U8081 ( .A(n5833), .Y(n3512) );
  BUFX2 U8082 ( .A(n5833), .Y(n3509) );
  BUFX2 U8083 ( .A(n5833), .Y(n3508) );
  BUFX2 U8084 ( .A(n5833), .Y(n3507) );
  BUFX2 U8085 ( .A(n5791), .Y(n3513) );
  BUFX2 U8086 ( .A(n5791), .Y(n3514) );
  BUFX2 U8087 ( .A(n5791), .Y(n3515) );
  BUFX2 U8088 ( .A(n5791), .Y(n3518) );
  BUFX2 U8089 ( .A(n5749), .Y(n3524) );
  BUFX2 U8090 ( .A(n5749), .Y(n3521) );
  BUFX2 U8091 ( .A(n5749), .Y(n3520) );
  BUFX2 U8092 ( .A(n5749), .Y(n3519) );
  BUFX2 U8093 ( .A(n5706), .Y(n3525) );
  BUFX2 U8094 ( .A(n5706), .Y(n3526) );
  BUFX2 U8095 ( .A(n5706), .Y(n3527) );
  BUFX2 U8096 ( .A(n5706), .Y(n3530) );
  BUFX2 U8097 ( .A(n6853), .Y(n3368) );
  BUFX2 U8098 ( .A(n6853), .Y(n3365) );
  BUFX2 U8099 ( .A(n6853), .Y(n3364) );
  BUFX2 U8100 ( .A(n6853), .Y(n3363) );
  BUFX2 U8101 ( .A(n6811), .Y(n3369) );
  BUFX2 U8102 ( .A(n6811), .Y(n3370) );
  BUFX2 U8103 ( .A(n6811), .Y(n3371) );
  BUFX2 U8104 ( .A(n6811), .Y(n3374) );
  BUFX2 U8105 ( .A(n6769), .Y(n3380) );
  BUFX2 U8106 ( .A(n6769), .Y(n3377) );
  BUFX2 U8107 ( .A(n6769), .Y(n3376) );
  BUFX2 U8108 ( .A(n6769), .Y(n3375) );
  BUFX2 U8109 ( .A(n6726), .Y(n3381) );
  BUFX2 U8110 ( .A(n6726), .Y(n3382) );
  BUFX2 U8111 ( .A(n6726), .Y(n3383) );
  BUFX2 U8112 ( .A(n6726), .Y(n3386) );
  BUFX2 U8113 ( .A(n6684), .Y(n3392) );
  BUFX2 U8114 ( .A(n6684), .Y(n3389) );
  BUFX2 U8115 ( .A(n6684), .Y(n3388) );
  BUFX2 U8116 ( .A(n6684), .Y(n3387) );
  BUFX2 U8117 ( .A(n6642), .Y(n3393) );
  BUFX2 U8118 ( .A(n6642), .Y(n3394) );
  BUFX2 U8119 ( .A(n6642), .Y(n3395) );
  BUFX2 U8120 ( .A(n6642), .Y(n3398) );
  BUFX2 U8121 ( .A(n6600), .Y(n3404) );
  BUFX2 U8122 ( .A(n6600), .Y(n3401) );
  BUFX2 U8123 ( .A(n6600), .Y(n3400) );
  BUFX2 U8124 ( .A(n6600), .Y(n3399) );
  BUFX2 U8125 ( .A(n6557), .Y(n3405) );
  BUFX2 U8126 ( .A(n6557), .Y(n3406) );
  BUFX2 U8127 ( .A(n6557), .Y(n3407) );
  BUFX2 U8128 ( .A(n6557), .Y(n3410) );
  BUFX2 U8129 ( .A(n6515), .Y(n3416) );
  BUFX2 U8130 ( .A(n6515), .Y(n3413) );
  BUFX2 U8131 ( .A(n6515), .Y(n3412) );
  BUFX2 U8132 ( .A(n6515), .Y(n3411) );
  BUFX2 U8133 ( .A(n6473), .Y(n3417) );
  BUFX2 U8134 ( .A(n6473), .Y(n3418) );
  BUFX2 U8135 ( .A(n6473), .Y(n3419) );
  BUFX2 U8136 ( .A(n6473), .Y(n3422) );
  BUFX2 U8137 ( .A(n6431), .Y(n3428) );
  BUFX2 U8138 ( .A(n6431), .Y(n3425) );
  BUFX2 U8139 ( .A(n6431), .Y(n3424) );
  BUFX2 U8140 ( .A(n6431), .Y(n3423) );
  BUFX2 U8141 ( .A(n6388), .Y(n3429) );
  BUFX2 U8142 ( .A(n6388), .Y(n3430) );
  BUFX2 U8143 ( .A(n6388), .Y(n3431) );
  BUFX2 U8144 ( .A(n6388), .Y(n3434) );
  BUFX2 U8145 ( .A(n6345), .Y(n3440) );
  BUFX2 U8146 ( .A(n6345), .Y(n3437) );
  BUFX2 U8147 ( .A(n6345), .Y(n3436) );
  BUFX2 U8148 ( .A(n6345), .Y(n3435) );
  BUFX2 U8149 ( .A(n6303), .Y(n3441) );
  BUFX2 U8150 ( .A(n6303), .Y(n3442) );
  BUFX2 U8151 ( .A(n6303), .Y(n3443) );
  BUFX2 U8152 ( .A(n6303), .Y(n3446) );
  BUFX2 U8153 ( .A(n6261), .Y(n3452) );
  BUFX2 U8154 ( .A(n6261), .Y(n3449) );
  BUFX2 U8155 ( .A(n6261), .Y(n3448) );
  BUFX2 U8156 ( .A(n6261), .Y(n3447) );
  BUFX2 U8157 ( .A(n6218), .Y(n3453) );
  BUFX2 U8158 ( .A(n6218), .Y(n3454) );
  BUFX2 U8159 ( .A(n6218), .Y(n3455) );
  BUFX2 U8160 ( .A(n6218), .Y(n3458) );
  AND2X2 U8161 ( .A(n5704), .B(n5705), .Y(n5574) );
  BUFX2 U8162 ( .A(n6940), .Y(n3356) );
  BUFX2 U8163 ( .A(n6897), .Y(n3362) );
  BUFX2 U8164 ( .A(n6897), .Y(n3358) );
  BUFX2 U8165 ( .A(n6897), .Y(n3359) );
  BUFX2 U8166 ( .A(n7532), .Y(n3267) );
  BUFX2 U8167 ( .A(n7532), .Y(n3268) );
  BUFX2 U8168 ( .A(n7532), .Y(n3269) );
  BUFX2 U8169 ( .A(n7532), .Y(n3272) );
  BUFX2 U8170 ( .A(n7490), .Y(n3278) );
  BUFX2 U8171 ( .A(n7490), .Y(n3275) );
  BUFX2 U8172 ( .A(n7490), .Y(n3274) );
  BUFX2 U8173 ( .A(n7490), .Y(n3273) );
  BUFX2 U8174 ( .A(n7448), .Y(n3279) );
  BUFX2 U8175 ( .A(n7448), .Y(n3280) );
  BUFX2 U8176 ( .A(n7448), .Y(n3281) );
  BUFX2 U8177 ( .A(n7448), .Y(n3284) );
  BUFX2 U8178 ( .A(n7405), .Y(n3290) );
  BUFX2 U8179 ( .A(n7405), .Y(n3287) );
  BUFX2 U8180 ( .A(n7405), .Y(n3286) );
  BUFX2 U8181 ( .A(n7405), .Y(n3285) );
  BUFX2 U8182 ( .A(n7363), .Y(n3291) );
  BUFX2 U8183 ( .A(n7363), .Y(n3292) );
  BUFX2 U8184 ( .A(n7363), .Y(n3293) );
  BUFX2 U8185 ( .A(n7363), .Y(n3296) );
  BUFX2 U8186 ( .A(n7321), .Y(n3302) );
  BUFX2 U8187 ( .A(n7321), .Y(n3299) );
  BUFX2 U8188 ( .A(n7321), .Y(n3298) );
  BUFX2 U8189 ( .A(n7321), .Y(n3297) );
  BUFX2 U8190 ( .A(n7279), .Y(n3303) );
  BUFX2 U8191 ( .A(n7279), .Y(n3304) );
  BUFX2 U8192 ( .A(n7279), .Y(n3305) );
  BUFX2 U8193 ( .A(n7279), .Y(n3308) );
  BUFX2 U8194 ( .A(n7236), .Y(n3314) );
  BUFX2 U8195 ( .A(n7236), .Y(n3311) );
  BUFX2 U8196 ( .A(n7236), .Y(n3310) );
  BUFX2 U8197 ( .A(n7236), .Y(n3309) );
  BUFX2 U8198 ( .A(n7194), .Y(n3315) );
  BUFX2 U8199 ( .A(n7194), .Y(n3316) );
  BUFX2 U8200 ( .A(n7194), .Y(n3317) );
  BUFX2 U8201 ( .A(n7194), .Y(n3320) );
  BUFX2 U8202 ( .A(n7152), .Y(n3326) );
  BUFX2 U8203 ( .A(n7152), .Y(n3323) );
  BUFX2 U8204 ( .A(n7152), .Y(n3322) );
  BUFX2 U8205 ( .A(n7152), .Y(n3321) );
  BUFX2 U8206 ( .A(n7110), .Y(n3327) );
  BUFX2 U8207 ( .A(n7110), .Y(n3328) );
  BUFX2 U8208 ( .A(n7110), .Y(n3329) );
  BUFX2 U8209 ( .A(n7110), .Y(n3332) );
  BUFX2 U8210 ( .A(n7067), .Y(n3338) );
  BUFX2 U8211 ( .A(n7067), .Y(n3335) );
  BUFX2 U8212 ( .A(n7067), .Y(n3334) );
  BUFX2 U8213 ( .A(n7067), .Y(n3333) );
  BUFX2 U8214 ( .A(n7024), .Y(n3339) );
  BUFX2 U8215 ( .A(n7024), .Y(n3340) );
  BUFX2 U8216 ( .A(n7024), .Y(n3341) );
  BUFX2 U8217 ( .A(n7024), .Y(n3344) );
  BUFX2 U8218 ( .A(n6982), .Y(n3350) );
  BUFX2 U8219 ( .A(n6982), .Y(n3347) );
  BUFX2 U8220 ( .A(n6982), .Y(n3346) );
  BUFX2 U8221 ( .A(n6982), .Y(n3345) );
  BUFX2 U8222 ( .A(n6940), .Y(n3351) );
  BUFX2 U8223 ( .A(n6897), .Y(n3357) );
  AND2X2 U8224 ( .A(wr_ptr[5]), .B(n6895), .Y(n7574) );
  BUFX2 U8225 ( .A(n8214), .Y(n3190) );
  BUFX2 U8226 ( .A(n8214), .Y(n3187) );
  BUFX2 U8227 ( .A(n8171), .Y(n3194) );
  BUFX2 U8228 ( .A(n8171), .Y(n3191) );
  BUFX2 U8229 ( .A(n8128), .Y(n3198) );
  BUFX2 U8230 ( .A(n8128), .Y(n3195) );
  BUFX2 U8231 ( .A(n8042), .Y(n3206) );
  BUFX2 U8232 ( .A(n8042), .Y(n3203) );
  BUFX2 U8233 ( .A(n8000), .Y(n3210) );
  BUFX2 U8234 ( .A(n8000), .Y(n3207) );
  BUFX2 U8235 ( .A(n7958), .Y(n3214) );
  BUFX2 U8236 ( .A(n7958), .Y(n3211) );
  BUFX2 U8237 ( .A(n7915), .Y(n3218) );
  BUFX2 U8238 ( .A(n7915), .Y(n3215) );
  BUFX2 U8239 ( .A(n7872), .Y(n3224) );
  BUFX2 U8240 ( .A(n7872), .Y(n3219) );
  BUFX2 U8241 ( .A(n7872), .Y(n3220) );
  BUFX2 U8242 ( .A(n7872), .Y(n3221) );
  BUFX2 U8243 ( .A(n7830), .Y(n3230) );
  BUFX2 U8244 ( .A(n7830), .Y(n3226) );
  BUFX2 U8245 ( .A(n7830), .Y(n3227) );
  BUFX2 U8246 ( .A(n7830), .Y(n3225) );
  BUFX2 U8247 ( .A(n7788), .Y(n3236) );
  BUFX2 U8248 ( .A(n7788), .Y(n3231) );
  BUFX2 U8249 ( .A(n7788), .Y(n3232) );
  BUFX2 U8250 ( .A(n7788), .Y(n3233) );
  BUFX2 U8251 ( .A(n7745), .Y(n3242) );
  BUFX2 U8252 ( .A(n7745), .Y(n3238) );
  BUFX2 U8253 ( .A(n7745), .Y(n3239) );
  BUFX2 U8254 ( .A(n7745), .Y(n3237) );
  BUFX2 U8255 ( .A(n7702), .Y(n3248) );
  BUFX2 U8256 ( .A(n7702), .Y(n3243) );
  BUFX2 U8257 ( .A(n7702), .Y(n3244) );
  BUFX2 U8258 ( .A(n7702), .Y(n3245) );
  BUFX2 U8259 ( .A(n7660), .Y(n3254) );
  BUFX2 U8260 ( .A(n7660), .Y(n3250) );
  BUFX2 U8261 ( .A(n7660), .Y(n3251) );
  BUFX2 U8262 ( .A(n7660), .Y(n3249) );
  BUFX2 U8263 ( .A(n7618), .Y(n3260) );
  BUFX2 U8264 ( .A(n7618), .Y(n3255) );
  BUFX2 U8265 ( .A(n7618), .Y(n3256) );
  BUFX2 U8266 ( .A(n7618), .Y(n3257) );
  AND2X2 U8267 ( .A(n6387), .B(n6215), .Y(n6768) );
  AND2X2 U8268 ( .A(n6387), .B(n6045), .Y(n6599) );
  AND2X2 U8269 ( .A(n6387), .B(n5875), .Y(n6430) );
  AND2X2 U8270 ( .A(n6387), .B(n5705), .Y(n6260) );
  AND2X2 U8271 ( .A(n6215), .B(n5704), .Y(n6088) );
  AND2X2 U8272 ( .A(n6045), .B(n5704), .Y(n5918) );
  AND2X2 U8273 ( .A(n5875), .B(n5704), .Y(n5748) );
  AND2X2 U8274 ( .A(n7066), .B(n6215), .Y(n7447) );
  AND2X2 U8275 ( .A(n7066), .B(n6045), .Y(n7278) );
  AND2X2 U8276 ( .A(n7066), .B(n5875), .Y(n7109) );
  AND2X2 U8277 ( .A(n7066), .B(n5705), .Y(n6939) );
  AND2X2 U8278 ( .A(n7744), .B(n6215), .Y(n8127) );
  INVX1 U8279 ( .A(fillcount[6]), .Y(n8277) );
  BUFX2 U8280 ( .A(n8085), .Y(n3202) );
  BUFX2 U8281 ( .A(n8085), .Y(n3199) );
  AND2X2 U8282 ( .A(n7744), .B(n6045), .Y(n7957) );
  AND2X2 U8283 ( .A(n7744), .B(n5875), .Y(n7787) );
  AND2X2 U8284 ( .A(n7744), .B(n5705), .Y(n7617) );
  INVX1 U8285 ( .A(fillcount[5]), .Y(n8267) );
  BUFX2 U8286 ( .A(n7575), .Y(n3266) );
  BUFX2 U8287 ( .A(n7575), .Y(n3261) );
  BUFX2 U8288 ( .A(n7575), .Y(n3262) );
  BUFX2 U8289 ( .A(n7575), .Y(n3263) );
  INVX4 U8290 ( .A(data_in[40]), .Y(n5571) );
  INVX4 U8291 ( .A(data_in[39]), .Y(n5569) );
  BUFX4 U8292 ( .A(n7872), .Y(n3222) );
  BUFX4 U8293 ( .A(n7872), .Y(n3223) );
  BUFX4 U8294 ( .A(n7830), .Y(n3228) );
  BUFX4 U8295 ( .A(n7830), .Y(n3229) );
  BUFX4 U8296 ( .A(n7788), .Y(n3234) );
  BUFX4 U8297 ( .A(n7788), .Y(n3235) );
  BUFX4 U8298 ( .A(n7745), .Y(n3240) );
  BUFX4 U8299 ( .A(n7745), .Y(n3241) );
  BUFX4 U8300 ( .A(n7702), .Y(n3246) );
  BUFX4 U8301 ( .A(n7702), .Y(n3247) );
  BUFX4 U8302 ( .A(n7660), .Y(n3252) );
  BUFX4 U8303 ( .A(n7660), .Y(n3253) );
  BUFX4 U8304 ( .A(n7618), .Y(n3258) );
  BUFX4 U8305 ( .A(n7618), .Y(n3259) );
  BUFX4 U8306 ( .A(n7575), .Y(n3264) );
  BUFX4 U8307 ( .A(n7575), .Y(n3265) );
  BUFX4 U8308 ( .A(n7532), .Y(n3270) );
  BUFX4 U8309 ( .A(n7532), .Y(n3271) );
  BUFX4 U8310 ( .A(n7490), .Y(n3276) );
  BUFX4 U8311 ( .A(n7490), .Y(n3277) );
  BUFX4 U8312 ( .A(n7448), .Y(n3282) );
  BUFX4 U8313 ( .A(n7448), .Y(n3283) );
  BUFX4 U8314 ( .A(n7405), .Y(n3288) );
  BUFX4 U8315 ( .A(n7405), .Y(n3289) );
  BUFX4 U8316 ( .A(n7363), .Y(n3294) );
  BUFX4 U8317 ( .A(n7363), .Y(n3295) );
  BUFX4 U8318 ( .A(n7321), .Y(n3300) );
  BUFX4 U8319 ( .A(n7321), .Y(n3301) );
  BUFX4 U8320 ( .A(n7279), .Y(n3306) );
  BUFX4 U8321 ( .A(n7279), .Y(n3307) );
  BUFX4 U8322 ( .A(n7236), .Y(n3312) );
  BUFX4 U8323 ( .A(n7236), .Y(n3313) );
  BUFX4 U8324 ( .A(n7194), .Y(n3318) );
  BUFX4 U8325 ( .A(n7194), .Y(n3319) );
  BUFX4 U8326 ( .A(n7152), .Y(n3324) );
  BUFX4 U8327 ( .A(n7152), .Y(n3325) );
  BUFX4 U8328 ( .A(n7110), .Y(n3330) );
  BUFX4 U8329 ( .A(n7110), .Y(n3331) );
  BUFX4 U8330 ( .A(n7067), .Y(n3336) );
  BUFX4 U8331 ( .A(n7067), .Y(n3337) );
  BUFX4 U8332 ( .A(n7024), .Y(n3342) );
  BUFX4 U8333 ( .A(n7024), .Y(n3343) );
  BUFX4 U8334 ( .A(n6982), .Y(n3348) );
  BUFX4 U8335 ( .A(n6982), .Y(n3349) );
  BUFX4 U8336 ( .A(n6940), .Y(n3354) );
  BUFX4 U8337 ( .A(n6940), .Y(n3355) );
  BUFX4 U8338 ( .A(n6897), .Y(n3360) );
  BUFX4 U8339 ( .A(n6897), .Y(n3361) );
  BUFX4 U8340 ( .A(n6853), .Y(n3366) );
  BUFX4 U8341 ( .A(n6853), .Y(n3367) );
  BUFX4 U8342 ( .A(n6811), .Y(n3372) );
  BUFX4 U8343 ( .A(n6811), .Y(n3373) );
  BUFX4 U8344 ( .A(n6769), .Y(n3378) );
  BUFX4 U8345 ( .A(n6769), .Y(n3379) );
  BUFX4 U8346 ( .A(n6726), .Y(n3384) );
  BUFX4 U8347 ( .A(n6726), .Y(n3385) );
  BUFX4 U8348 ( .A(n6684), .Y(n3390) );
  BUFX4 U8349 ( .A(n6684), .Y(n3391) );
  BUFX4 U8350 ( .A(n6642), .Y(n3396) );
  BUFX4 U8351 ( .A(n6642), .Y(n3397) );
  BUFX4 U8352 ( .A(n6600), .Y(n3402) );
  BUFX4 U8353 ( .A(n6600), .Y(n3403) );
  BUFX4 U8354 ( .A(n6557), .Y(n3408) );
  BUFX4 U8355 ( .A(n6557), .Y(n3409) );
  BUFX4 U8356 ( .A(n6515), .Y(n3414) );
  BUFX4 U8357 ( .A(n6515), .Y(n3415) );
  BUFX4 U8358 ( .A(n6473), .Y(n3420) );
  BUFX4 U8359 ( .A(n6473), .Y(n3421) );
  BUFX4 U8360 ( .A(n6431), .Y(n3426) );
  BUFX4 U8361 ( .A(n6431), .Y(n3427) );
  BUFX4 U8362 ( .A(n6388), .Y(n3432) );
  BUFX4 U8363 ( .A(n6388), .Y(n3433) );
  BUFX4 U8364 ( .A(n6345), .Y(n3438) );
  BUFX4 U8365 ( .A(n6345), .Y(n3439) );
  BUFX4 U8366 ( .A(n6303), .Y(n3444) );
  BUFX4 U8367 ( .A(n6303), .Y(n3445) );
  BUFX4 U8368 ( .A(n6261), .Y(n3450) );
  BUFX4 U8369 ( .A(n6261), .Y(n3451) );
  BUFX4 U8370 ( .A(n6218), .Y(n3456) );
  BUFX4 U8371 ( .A(n6218), .Y(n3457) );
  BUFX4 U8372 ( .A(n6173), .Y(n3462) );
  BUFX4 U8373 ( .A(n6173), .Y(n3463) );
  BUFX4 U8374 ( .A(n6131), .Y(n3468) );
  BUFX4 U8375 ( .A(n6131), .Y(n3469) );
  BUFX4 U8376 ( .A(n6089), .Y(n3474) );
  BUFX4 U8377 ( .A(n6089), .Y(n3475) );
  BUFX4 U8378 ( .A(n6046), .Y(n3480) );
  BUFX4 U8379 ( .A(n6046), .Y(n3481) );
  BUFX4 U8380 ( .A(n6003), .Y(n3486) );
  BUFX4 U8381 ( .A(n6003), .Y(n3487) );
  BUFX4 U8382 ( .A(n5961), .Y(n3492) );
  BUFX4 U8383 ( .A(n5961), .Y(n3493) );
  BUFX4 U8384 ( .A(n5919), .Y(n3498) );
  BUFX4 U8385 ( .A(n5919), .Y(n3499) );
  BUFX4 U8386 ( .A(n5876), .Y(n3504) );
  BUFX4 U8387 ( .A(n5876), .Y(n3505) );
  BUFX4 U8388 ( .A(n5833), .Y(n3510) );
  BUFX4 U8389 ( .A(n5833), .Y(n3511) );
  BUFX4 U8390 ( .A(n5791), .Y(n3516) );
  BUFX4 U8391 ( .A(n5791), .Y(n3517) );
  BUFX4 U8392 ( .A(n5749), .Y(n3522) );
  BUFX4 U8393 ( .A(n5749), .Y(n3523) );
  BUFX4 U8394 ( .A(n5706), .Y(n3528) );
  BUFX4 U8395 ( .A(n5706), .Y(n3529) );
  BUFX4 U8396 ( .A(n5661), .Y(n3534) );
  BUFX4 U8397 ( .A(n5661), .Y(n3535) );
  BUFX4 U8398 ( .A(n5618), .Y(n3540) );
  BUFX4 U8399 ( .A(n5618), .Y(n3541) );
  BUFX4 U8400 ( .A(n5575), .Y(n3546) );
  BUFX4 U8401 ( .A(n5575), .Y(n3547) );
  BUFX4 U8402 ( .A(n5490), .Y(n3552) );
  BUFX4 U8403 ( .A(n5490), .Y(n3553) );
endmodule


module FIFO_DEPTH_P26_WIDTH33 ( clk, reset, data_in, put, get, data_out, empty, 
        full, fillcount );
  input [32:0] data_in;
  output [32:0] data_out;
  output [6:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   n13, n14, n15, n16, n17, n18, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6504, n6573, n6642, n6677, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816;
  wire   [5:0] wr_ptr;
  wire   [2111:0] arr;

  DFFPOSX1 fillcount_reg_0_ ( .D(n8882), .CLK(clk), .Q(fillcount[0]) );
  DFFPOSX1 fillcount_reg_1_ ( .D(n8881), .CLK(clk), .Q(fillcount[1]) );
  DFFPOSX1 fillcount_reg_6_ ( .D(n8880), .CLK(clk), .Q(fillcount[6]) );
  DFFPOSX1 fillcount_reg_2_ ( .D(n8879), .CLK(clk), .Q(fillcount[2]) );
  DFFPOSX1 fillcount_reg_3_ ( .D(n8878), .CLK(clk), .Q(fillcount[3]) );
  DFFPOSX1 fillcount_reg_4_ ( .D(n8877), .CLK(clk), .Q(fillcount[4]) );
  DFFPOSX1 fillcount_reg_5_ ( .D(n8876), .CLK(clk), .Q(fillcount[5]) );
  DFFPOSX1 wr_ptr_reg_0_ ( .D(n8875), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n8874), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n8873), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n8872), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n8871), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 wr_ptr_reg_5_ ( .D(n8870), .CLK(clk), .Q(wr_ptr[5]) );
  DFFPOSX1 arr_reg_63__32_ ( .D(n219), .CLK(clk), .Q(arr[2111]) );
  DFFPOSX1 arr_reg_63__31_ ( .D(n347), .CLK(clk), .Q(arr[2110]) );
  DFFPOSX1 arr_reg_63__30_ ( .D(n346), .CLK(clk), .Q(arr[2109]) );
  DFFPOSX1 arr_reg_63__29_ ( .D(n345), .CLK(clk), .Q(arr[2108]) );
  DFFPOSX1 arr_reg_63__28_ ( .D(n344), .CLK(clk), .Q(arr[2107]) );
  DFFPOSX1 arr_reg_63__27_ ( .D(n343), .CLK(clk), .Q(arr[2106]) );
  DFFPOSX1 arr_reg_63__26_ ( .D(n342), .CLK(clk), .Q(arr[2105]) );
  DFFPOSX1 arr_reg_63__25_ ( .D(n341), .CLK(clk), .Q(arr[2104]) );
  DFFPOSX1 arr_reg_63__24_ ( .D(n340), .CLK(clk), .Q(arr[2103]) );
  DFFPOSX1 arr_reg_63__23_ ( .D(n339), .CLK(clk), .Q(arr[2102]) );
  DFFPOSX1 arr_reg_63__22_ ( .D(n218), .CLK(clk), .Q(arr[2101]) );
  DFFPOSX1 arr_reg_63__21_ ( .D(n217), .CLK(clk), .Q(arr[2100]) );
  DFFPOSX1 arr_reg_63__20_ ( .D(n216), .CLK(clk), .Q(arr[2099]) );
  DFFPOSX1 arr_reg_63__19_ ( .D(n215), .CLK(clk), .Q(arr[2098]) );
  DFFPOSX1 arr_reg_63__18_ ( .D(n214), .CLK(clk), .Q(arr[2097]) );
  DFFPOSX1 arr_reg_63__17_ ( .D(n213), .CLK(clk), .Q(arr[2096]) );
  DFFPOSX1 arr_reg_63__16_ ( .D(n212), .CLK(clk), .Q(arr[2095]) );
  DFFPOSX1 arr_reg_63__15_ ( .D(n211), .CLK(clk), .Q(arr[2094]) );
  DFFPOSX1 arr_reg_63__14_ ( .D(n210), .CLK(clk), .Q(arr[2093]) );
  DFFPOSX1 arr_reg_63__13_ ( .D(n209), .CLK(clk), .Q(arr[2092]) );
  DFFPOSX1 arr_reg_63__12_ ( .D(n208), .CLK(clk), .Q(arr[2091]) );
  DFFPOSX1 arr_reg_63__11_ ( .D(n207), .CLK(clk), .Q(arr[2090]) );
  DFFPOSX1 arr_reg_63__10_ ( .D(n206), .CLK(clk), .Q(arr[2089]) );
  DFFPOSX1 arr_reg_63__9_ ( .D(n205), .CLK(clk), .Q(arr[2088]) );
  DFFPOSX1 arr_reg_63__8_ ( .D(n338), .CLK(clk), .Q(arr[2087]) );
  DFFPOSX1 arr_reg_63__7_ ( .D(n337), .CLK(clk), .Q(arr[2086]) );
  DFFPOSX1 arr_reg_63__6_ ( .D(n204), .CLK(clk), .Q(arr[2085]) );
  DFFPOSX1 arr_reg_63__5_ ( .D(n203), .CLK(clk), .Q(arr[2084]) );
  DFFPOSX1 arr_reg_63__4_ ( .D(n336), .CLK(clk), .Q(arr[2083]) );
  DFFPOSX1 arr_reg_63__3_ ( .D(n335), .CLK(clk), .Q(arr[2082]) );
  DFFPOSX1 arr_reg_63__2_ ( .D(n334), .CLK(clk), .Q(arr[2081]) );
  DFFPOSX1 arr_reg_63__1_ ( .D(n333), .CLK(clk), .Q(arr[2080]) );
  DFFPOSX1 arr_reg_63__0_ ( .D(n332), .CLK(clk), .Q(arr[2079]) );
  DFFPOSX1 arr_reg_62__32_ ( .D(n202), .CLK(clk), .Q(arr[2078]) );
  DFFPOSX1 arr_reg_62__31_ ( .D(n331), .CLK(clk), .Q(arr[2077]) );
  DFFPOSX1 arr_reg_62__30_ ( .D(n330), .CLK(clk), .Q(arr[2076]) );
  DFFPOSX1 arr_reg_62__29_ ( .D(n329), .CLK(clk), .Q(arr[2075]) );
  DFFPOSX1 arr_reg_62__28_ ( .D(n328), .CLK(clk), .Q(arr[2074]) );
  DFFPOSX1 arr_reg_62__27_ ( .D(n327), .CLK(clk), .Q(arr[2073]) );
  DFFPOSX1 arr_reg_62__26_ ( .D(n326), .CLK(clk), .Q(arr[2072]) );
  DFFPOSX1 arr_reg_62__25_ ( .D(n325), .CLK(clk), .Q(arr[2071]) );
  DFFPOSX1 arr_reg_62__24_ ( .D(n324), .CLK(clk), .Q(arr[2070]) );
  DFFPOSX1 arr_reg_62__23_ ( .D(n323), .CLK(clk), .Q(arr[2069]) );
  DFFPOSX1 arr_reg_62__22_ ( .D(n201), .CLK(clk), .Q(arr[2068]) );
  DFFPOSX1 arr_reg_62__21_ ( .D(n200), .CLK(clk), .Q(arr[2067]) );
  DFFPOSX1 arr_reg_62__20_ ( .D(n199), .CLK(clk), .Q(arr[2066]) );
  DFFPOSX1 arr_reg_62__19_ ( .D(n198), .CLK(clk), .Q(arr[2065]) );
  DFFPOSX1 arr_reg_62__18_ ( .D(n197), .CLK(clk), .Q(arr[2064]) );
  DFFPOSX1 arr_reg_62__17_ ( .D(n196), .CLK(clk), .Q(arr[2063]) );
  DFFPOSX1 arr_reg_62__16_ ( .D(n195), .CLK(clk), .Q(arr[2062]) );
  DFFPOSX1 arr_reg_62__15_ ( .D(n194), .CLK(clk), .Q(arr[2061]) );
  DFFPOSX1 arr_reg_62__14_ ( .D(n193), .CLK(clk), .Q(arr[2060]) );
  DFFPOSX1 arr_reg_62__13_ ( .D(n192), .CLK(clk), .Q(arr[2059]) );
  DFFPOSX1 arr_reg_62__12_ ( .D(n191), .CLK(clk), .Q(arr[2058]) );
  DFFPOSX1 arr_reg_62__11_ ( .D(n190), .CLK(clk), .Q(arr[2057]) );
  DFFPOSX1 arr_reg_62__10_ ( .D(n189), .CLK(clk), .Q(arr[2056]) );
  DFFPOSX1 arr_reg_62__9_ ( .D(n188), .CLK(clk), .Q(arr[2055]) );
  DFFPOSX1 arr_reg_62__8_ ( .D(n322), .CLK(clk), .Q(arr[2054]) );
  DFFPOSX1 arr_reg_62__7_ ( .D(n321), .CLK(clk), .Q(arr[2053]) );
  DFFPOSX1 arr_reg_62__6_ ( .D(n187), .CLK(clk), .Q(arr[2052]) );
  DFFPOSX1 arr_reg_62__5_ ( .D(n186), .CLK(clk), .Q(arr[2051]) );
  DFFPOSX1 arr_reg_62__4_ ( .D(n320), .CLK(clk), .Q(arr[2050]) );
  DFFPOSX1 arr_reg_62__3_ ( .D(n319), .CLK(clk), .Q(arr[2049]) );
  DFFPOSX1 arr_reg_62__2_ ( .D(n318), .CLK(clk), .Q(arr[2048]) );
  DFFPOSX1 arr_reg_62__1_ ( .D(n317), .CLK(clk), .Q(arr[2047]) );
  DFFPOSX1 arr_reg_62__0_ ( .D(n316), .CLK(clk), .Q(arr[2046]) );
  DFFPOSX1 arr_reg_61__32_ ( .D(n185), .CLK(clk), .Q(arr[2045]) );
  DFFPOSX1 arr_reg_61__31_ ( .D(n315), .CLK(clk), .Q(arr[2044]) );
  DFFPOSX1 arr_reg_61__30_ ( .D(n314), .CLK(clk), .Q(arr[2043]) );
  DFFPOSX1 arr_reg_61__29_ ( .D(n313), .CLK(clk), .Q(arr[2042]) );
  DFFPOSX1 arr_reg_61__28_ ( .D(n312), .CLK(clk), .Q(arr[2041]) );
  DFFPOSX1 arr_reg_61__27_ ( .D(n311), .CLK(clk), .Q(arr[2040]) );
  DFFPOSX1 arr_reg_61__26_ ( .D(n310), .CLK(clk), .Q(arr[2039]) );
  DFFPOSX1 arr_reg_61__25_ ( .D(n309), .CLK(clk), .Q(arr[2038]) );
  DFFPOSX1 arr_reg_61__24_ ( .D(n308), .CLK(clk), .Q(arr[2037]) );
  DFFPOSX1 arr_reg_61__23_ ( .D(n307), .CLK(clk), .Q(arr[2036]) );
  DFFPOSX1 arr_reg_61__22_ ( .D(n184), .CLK(clk), .Q(arr[2035]) );
  DFFPOSX1 arr_reg_61__21_ ( .D(n183), .CLK(clk), .Q(arr[2034]) );
  DFFPOSX1 arr_reg_61__20_ ( .D(n182), .CLK(clk), .Q(arr[2033]) );
  DFFPOSX1 arr_reg_61__19_ ( .D(n181), .CLK(clk), .Q(arr[2032]) );
  DFFPOSX1 arr_reg_61__18_ ( .D(n180), .CLK(clk), .Q(arr[2031]) );
  DFFPOSX1 arr_reg_61__17_ ( .D(n179), .CLK(clk), .Q(arr[2030]) );
  DFFPOSX1 arr_reg_61__16_ ( .D(n178), .CLK(clk), .Q(arr[2029]) );
  DFFPOSX1 arr_reg_61__15_ ( .D(n177), .CLK(clk), .Q(arr[2028]) );
  DFFPOSX1 arr_reg_61__14_ ( .D(n176), .CLK(clk), .Q(arr[2027]) );
  DFFPOSX1 arr_reg_61__13_ ( .D(n175), .CLK(clk), .Q(arr[2026]) );
  DFFPOSX1 arr_reg_61__12_ ( .D(n174), .CLK(clk), .Q(arr[2025]) );
  DFFPOSX1 arr_reg_61__11_ ( .D(n173), .CLK(clk), .Q(arr[2024]) );
  DFFPOSX1 arr_reg_61__10_ ( .D(n172), .CLK(clk), .Q(arr[2023]) );
  DFFPOSX1 arr_reg_61__9_ ( .D(n171), .CLK(clk), .Q(arr[2022]) );
  DFFPOSX1 arr_reg_61__8_ ( .D(n306), .CLK(clk), .Q(arr[2021]) );
  DFFPOSX1 arr_reg_61__7_ ( .D(n305), .CLK(clk), .Q(arr[2020]) );
  DFFPOSX1 arr_reg_61__6_ ( .D(n170), .CLK(clk), .Q(arr[2019]) );
  DFFPOSX1 arr_reg_61__5_ ( .D(n169), .CLK(clk), .Q(arr[2018]) );
  DFFPOSX1 arr_reg_61__4_ ( .D(n304), .CLK(clk), .Q(arr[2017]) );
  DFFPOSX1 arr_reg_61__3_ ( .D(n303), .CLK(clk), .Q(arr[2016]) );
  DFFPOSX1 arr_reg_61__2_ ( .D(n302), .CLK(clk), .Q(arr[2015]) );
  DFFPOSX1 arr_reg_61__1_ ( .D(n301), .CLK(clk), .Q(arr[2014]) );
  DFFPOSX1 arr_reg_61__0_ ( .D(n300), .CLK(clk), .Q(arr[2013]) );
  DFFPOSX1 arr_reg_60__32_ ( .D(n168), .CLK(clk), .Q(arr[2012]) );
  DFFPOSX1 arr_reg_60__31_ ( .D(n299), .CLK(clk), .Q(arr[2011]) );
  DFFPOSX1 arr_reg_60__30_ ( .D(n298), .CLK(clk), .Q(arr[2010]) );
  DFFPOSX1 arr_reg_60__29_ ( .D(n297), .CLK(clk), .Q(arr[2009]) );
  DFFPOSX1 arr_reg_60__28_ ( .D(n296), .CLK(clk), .Q(arr[2008]) );
  DFFPOSX1 arr_reg_60__27_ ( .D(n295), .CLK(clk), .Q(arr[2007]) );
  DFFPOSX1 arr_reg_60__26_ ( .D(n294), .CLK(clk), .Q(arr[2006]) );
  DFFPOSX1 arr_reg_60__25_ ( .D(n293), .CLK(clk), .Q(arr[2005]) );
  DFFPOSX1 arr_reg_60__24_ ( .D(n292), .CLK(clk), .Q(arr[2004]) );
  DFFPOSX1 arr_reg_60__23_ ( .D(n291), .CLK(clk), .Q(arr[2003]) );
  DFFPOSX1 arr_reg_60__22_ ( .D(n167), .CLK(clk), .Q(arr[2002]) );
  DFFPOSX1 arr_reg_60__21_ ( .D(n166), .CLK(clk), .Q(arr[2001]) );
  DFFPOSX1 arr_reg_60__20_ ( .D(n165), .CLK(clk), .Q(arr[2000]) );
  DFFPOSX1 arr_reg_60__19_ ( .D(n164), .CLK(clk), .Q(arr[1999]) );
  DFFPOSX1 arr_reg_60__18_ ( .D(n163), .CLK(clk), .Q(arr[1998]) );
  DFFPOSX1 arr_reg_60__17_ ( .D(n162), .CLK(clk), .Q(arr[1997]) );
  DFFPOSX1 arr_reg_60__16_ ( .D(n161), .CLK(clk), .Q(arr[1996]) );
  DFFPOSX1 arr_reg_60__15_ ( .D(n160), .CLK(clk), .Q(arr[1995]) );
  DFFPOSX1 arr_reg_60__14_ ( .D(n159), .CLK(clk), .Q(arr[1994]) );
  DFFPOSX1 arr_reg_60__13_ ( .D(n158), .CLK(clk), .Q(arr[1993]) );
  DFFPOSX1 arr_reg_60__12_ ( .D(n157), .CLK(clk), .Q(arr[1992]) );
  DFFPOSX1 arr_reg_60__11_ ( .D(n156), .CLK(clk), .Q(arr[1991]) );
  DFFPOSX1 arr_reg_60__10_ ( .D(n155), .CLK(clk), .Q(arr[1990]) );
  DFFPOSX1 arr_reg_60__9_ ( .D(n154), .CLK(clk), .Q(arr[1989]) );
  DFFPOSX1 arr_reg_60__8_ ( .D(n290), .CLK(clk), .Q(arr[1988]) );
  DFFPOSX1 arr_reg_60__7_ ( .D(n289), .CLK(clk), .Q(arr[1987]) );
  DFFPOSX1 arr_reg_60__6_ ( .D(n153), .CLK(clk), .Q(arr[1986]) );
  DFFPOSX1 arr_reg_60__5_ ( .D(n152), .CLK(clk), .Q(arr[1985]) );
  DFFPOSX1 arr_reg_60__4_ ( .D(n288), .CLK(clk), .Q(arr[1984]) );
  DFFPOSX1 arr_reg_60__3_ ( .D(n287), .CLK(clk), .Q(arr[1983]) );
  DFFPOSX1 arr_reg_60__2_ ( .D(n286), .CLK(clk), .Q(arr[1982]) );
  DFFPOSX1 arr_reg_60__1_ ( .D(n285), .CLK(clk), .Q(arr[1981]) );
  DFFPOSX1 arr_reg_60__0_ ( .D(n284), .CLK(clk), .Q(arr[1980]) );
  DFFPOSX1 arr_reg_59__32_ ( .D(n151), .CLK(clk), .Q(arr[1979]) );
  DFFPOSX1 arr_reg_59__31_ ( .D(n283), .CLK(clk), .Q(arr[1978]) );
  DFFPOSX1 arr_reg_59__30_ ( .D(n282), .CLK(clk), .Q(arr[1977]) );
  DFFPOSX1 arr_reg_59__29_ ( .D(n281), .CLK(clk), .Q(arr[1976]) );
  DFFPOSX1 arr_reg_59__28_ ( .D(n280), .CLK(clk), .Q(arr[1975]) );
  DFFPOSX1 arr_reg_59__27_ ( .D(n279), .CLK(clk), .Q(arr[1974]) );
  DFFPOSX1 arr_reg_59__26_ ( .D(n278), .CLK(clk), .Q(arr[1973]) );
  DFFPOSX1 arr_reg_59__25_ ( .D(n277), .CLK(clk), .Q(arr[1972]) );
  DFFPOSX1 arr_reg_59__24_ ( .D(n276), .CLK(clk), .Q(arr[1971]) );
  DFFPOSX1 arr_reg_59__23_ ( .D(n275), .CLK(clk), .Q(arr[1970]) );
  DFFPOSX1 arr_reg_59__22_ ( .D(n150), .CLK(clk), .Q(arr[1969]) );
  DFFPOSX1 arr_reg_59__21_ ( .D(n149), .CLK(clk), .Q(arr[1968]) );
  DFFPOSX1 arr_reg_59__20_ ( .D(n148), .CLK(clk), .Q(arr[1967]) );
  DFFPOSX1 arr_reg_59__19_ ( .D(n147), .CLK(clk), .Q(arr[1966]) );
  DFFPOSX1 arr_reg_59__18_ ( .D(n146), .CLK(clk), .Q(arr[1965]) );
  DFFPOSX1 arr_reg_59__17_ ( .D(n145), .CLK(clk), .Q(arr[1964]) );
  DFFPOSX1 arr_reg_59__16_ ( .D(n144), .CLK(clk), .Q(arr[1963]) );
  DFFPOSX1 arr_reg_59__15_ ( .D(n143), .CLK(clk), .Q(arr[1962]) );
  DFFPOSX1 arr_reg_59__14_ ( .D(n142), .CLK(clk), .Q(arr[1961]) );
  DFFPOSX1 arr_reg_59__13_ ( .D(n141), .CLK(clk), .Q(arr[1960]) );
  DFFPOSX1 arr_reg_59__12_ ( .D(n140), .CLK(clk), .Q(arr[1959]) );
  DFFPOSX1 arr_reg_59__11_ ( .D(n139), .CLK(clk), .Q(arr[1958]) );
  DFFPOSX1 arr_reg_59__10_ ( .D(n138), .CLK(clk), .Q(arr[1957]) );
  DFFPOSX1 arr_reg_59__9_ ( .D(n137), .CLK(clk), .Q(arr[1956]) );
  DFFPOSX1 arr_reg_59__8_ ( .D(n274), .CLK(clk), .Q(arr[1955]) );
  DFFPOSX1 arr_reg_59__7_ ( .D(n273), .CLK(clk), .Q(arr[1954]) );
  DFFPOSX1 arr_reg_59__6_ ( .D(n136), .CLK(clk), .Q(arr[1953]) );
  DFFPOSX1 arr_reg_59__5_ ( .D(n135), .CLK(clk), .Q(arr[1952]) );
  DFFPOSX1 arr_reg_59__4_ ( .D(n272), .CLK(clk), .Q(arr[1951]) );
  DFFPOSX1 arr_reg_59__3_ ( .D(n271), .CLK(clk), .Q(arr[1950]) );
  DFFPOSX1 arr_reg_59__2_ ( .D(n270), .CLK(clk), .Q(arr[1949]) );
  DFFPOSX1 arr_reg_59__1_ ( .D(n269), .CLK(clk), .Q(arr[1948]) );
  DFFPOSX1 arr_reg_59__0_ ( .D(n268), .CLK(clk), .Q(arr[1947]) );
  DFFPOSX1 arr_reg_58__32_ ( .D(n134), .CLK(clk), .Q(arr[1946]) );
  DFFPOSX1 arr_reg_58__31_ ( .D(n267), .CLK(clk), .Q(arr[1945]) );
  DFFPOSX1 arr_reg_58__30_ ( .D(n266), .CLK(clk), .Q(arr[1944]) );
  DFFPOSX1 arr_reg_58__29_ ( .D(n265), .CLK(clk), .Q(arr[1943]) );
  DFFPOSX1 arr_reg_58__28_ ( .D(n264), .CLK(clk), .Q(arr[1942]) );
  DFFPOSX1 arr_reg_58__27_ ( .D(n263), .CLK(clk), .Q(arr[1941]) );
  DFFPOSX1 arr_reg_58__26_ ( .D(n262), .CLK(clk), .Q(arr[1940]) );
  DFFPOSX1 arr_reg_58__25_ ( .D(n261), .CLK(clk), .Q(arr[1939]) );
  DFFPOSX1 arr_reg_58__24_ ( .D(n260), .CLK(clk), .Q(arr[1938]) );
  DFFPOSX1 arr_reg_58__23_ ( .D(n259), .CLK(clk), .Q(arr[1937]) );
  DFFPOSX1 arr_reg_58__22_ ( .D(n133), .CLK(clk), .Q(arr[1936]) );
  DFFPOSX1 arr_reg_58__21_ ( .D(n132), .CLK(clk), .Q(arr[1935]) );
  DFFPOSX1 arr_reg_58__20_ ( .D(n131), .CLK(clk), .Q(arr[1934]) );
  DFFPOSX1 arr_reg_58__19_ ( .D(n130), .CLK(clk), .Q(arr[1933]) );
  DFFPOSX1 arr_reg_58__18_ ( .D(n129), .CLK(clk), .Q(arr[1932]) );
  DFFPOSX1 arr_reg_58__17_ ( .D(n128), .CLK(clk), .Q(arr[1931]) );
  DFFPOSX1 arr_reg_58__16_ ( .D(n127), .CLK(clk), .Q(arr[1930]) );
  DFFPOSX1 arr_reg_58__15_ ( .D(n126), .CLK(clk), .Q(arr[1929]) );
  DFFPOSX1 arr_reg_58__14_ ( .D(n125), .CLK(clk), .Q(arr[1928]) );
  DFFPOSX1 arr_reg_58__13_ ( .D(n124), .CLK(clk), .Q(arr[1927]) );
  DFFPOSX1 arr_reg_58__12_ ( .D(n123), .CLK(clk), .Q(arr[1926]) );
  DFFPOSX1 arr_reg_58__11_ ( .D(n122), .CLK(clk), .Q(arr[1925]) );
  DFFPOSX1 arr_reg_58__10_ ( .D(n121), .CLK(clk), .Q(arr[1924]) );
  DFFPOSX1 arr_reg_58__9_ ( .D(n120), .CLK(clk), .Q(arr[1923]) );
  DFFPOSX1 arr_reg_58__8_ ( .D(n258), .CLK(clk), .Q(arr[1922]) );
  DFFPOSX1 arr_reg_58__7_ ( .D(n257), .CLK(clk), .Q(arr[1921]) );
  DFFPOSX1 arr_reg_58__6_ ( .D(n119), .CLK(clk), .Q(arr[1920]) );
  DFFPOSX1 arr_reg_58__5_ ( .D(n118), .CLK(clk), .Q(arr[1919]) );
  DFFPOSX1 arr_reg_58__4_ ( .D(n256), .CLK(clk), .Q(arr[1918]) );
  DFFPOSX1 arr_reg_58__3_ ( .D(n255), .CLK(clk), .Q(arr[1917]) );
  DFFPOSX1 arr_reg_58__2_ ( .D(n254), .CLK(clk), .Q(arr[1916]) );
  DFFPOSX1 arr_reg_58__1_ ( .D(n253), .CLK(clk), .Q(arr[1915]) );
  DFFPOSX1 arr_reg_58__0_ ( .D(n252), .CLK(clk), .Q(arr[1914]) );
  DFFPOSX1 arr_reg_57__32_ ( .D(n117), .CLK(clk), .Q(arr[1913]) );
  DFFPOSX1 arr_reg_57__31_ ( .D(n251), .CLK(clk), .Q(arr[1912]) );
  DFFPOSX1 arr_reg_57__30_ ( .D(n250), .CLK(clk), .Q(arr[1911]) );
  DFFPOSX1 arr_reg_57__29_ ( .D(n249), .CLK(clk), .Q(arr[1910]) );
  DFFPOSX1 arr_reg_57__28_ ( .D(n248), .CLK(clk), .Q(arr[1909]) );
  DFFPOSX1 arr_reg_57__27_ ( .D(n247), .CLK(clk), .Q(arr[1908]) );
  DFFPOSX1 arr_reg_57__26_ ( .D(n246), .CLK(clk), .Q(arr[1907]) );
  DFFPOSX1 arr_reg_57__25_ ( .D(n245), .CLK(clk), .Q(arr[1906]) );
  DFFPOSX1 arr_reg_57__24_ ( .D(n244), .CLK(clk), .Q(arr[1905]) );
  DFFPOSX1 arr_reg_57__23_ ( .D(n243), .CLK(clk), .Q(arr[1904]) );
  DFFPOSX1 arr_reg_57__22_ ( .D(n116), .CLK(clk), .Q(arr[1903]) );
  DFFPOSX1 arr_reg_57__21_ ( .D(n115), .CLK(clk), .Q(arr[1902]) );
  DFFPOSX1 arr_reg_57__20_ ( .D(n114), .CLK(clk), .Q(arr[1901]) );
  DFFPOSX1 arr_reg_57__19_ ( .D(n113), .CLK(clk), .Q(arr[1900]) );
  DFFPOSX1 arr_reg_57__18_ ( .D(n112), .CLK(clk), .Q(arr[1899]) );
  DFFPOSX1 arr_reg_57__17_ ( .D(n111), .CLK(clk), .Q(arr[1898]) );
  DFFPOSX1 arr_reg_57__16_ ( .D(n110), .CLK(clk), .Q(arr[1897]) );
  DFFPOSX1 arr_reg_57__15_ ( .D(n109), .CLK(clk), .Q(arr[1896]) );
  DFFPOSX1 arr_reg_57__14_ ( .D(n108), .CLK(clk), .Q(arr[1895]) );
  DFFPOSX1 arr_reg_57__13_ ( .D(n107), .CLK(clk), .Q(arr[1894]) );
  DFFPOSX1 arr_reg_57__12_ ( .D(n106), .CLK(clk), .Q(arr[1893]) );
  DFFPOSX1 arr_reg_57__11_ ( .D(n105), .CLK(clk), .Q(arr[1892]) );
  DFFPOSX1 arr_reg_57__10_ ( .D(n104), .CLK(clk), .Q(arr[1891]) );
  DFFPOSX1 arr_reg_57__9_ ( .D(n103), .CLK(clk), .Q(arr[1890]) );
  DFFPOSX1 arr_reg_57__8_ ( .D(n242), .CLK(clk), .Q(arr[1889]) );
  DFFPOSX1 arr_reg_57__7_ ( .D(n241), .CLK(clk), .Q(arr[1888]) );
  DFFPOSX1 arr_reg_57__6_ ( .D(n102), .CLK(clk), .Q(arr[1887]) );
  DFFPOSX1 arr_reg_57__5_ ( .D(n101), .CLK(clk), .Q(arr[1886]) );
  DFFPOSX1 arr_reg_57__4_ ( .D(n240), .CLK(clk), .Q(arr[1885]) );
  DFFPOSX1 arr_reg_57__3_ ( .D(n239), .CLK(clk), .Q(arr[1884]) );
  DFFPOSX1 arr_reg_57__2_ ( .D(n238), .CLK(clk), .Q(arr[1883]) );
  DFFPOSX1 arr_reg_57__1_ ( .D(n237), .CLK(clk), .Q(arr[1882]) );
  DFFPOSX1 arr_reg_57__0_ ( .D(n236), .CLK(clk), .Q(arr[1881]) );
  DFFPOSX1 arr_reg_56__32_ ( .D(n100), .CLK(clk), .Q(arr[1880]) );
  DFFPOSX1 arr_reg_56__31_ ( .D(n235), .CLK(clk), .Q(arr[1879]) );
  DFFPOSX1 arr_reg_56__30_ ( .D(n234), .CLK(clk), .Q(arr[1878]) );
  DFFPOSX1 arr_reg_56__29_ ( .D(n233), .CLK(clk), .Q(arr[1877]) );
  DFFPOSX1 arr_reg_56__28_ ( .D(n232), .CLK(clk), .Q(arr[1876]) );
  DFFPOSX1 arr_reg_56__27_ ( .D(n231), .CLK(clk), .Q(arr[1875]) );
  DFFPOSX1 arr_reg_56__26_ ( .D(n230), .CLK(clk), .Q(arr[1874]) );
  DFFPOSX1 arr_reg_56__25_ ( .D(n229), .CLK(clk), .Q(arr[1873]) );
  DFFPOSX1 arr_reg_56__24_ ( .D(n228), .CLK(clk), .Q(arr[1872]) );
  DFFPOSX1 arr_reg_56__23_ ( .D(n227), .CLK(clk), .Q(arr[1871]) );
  DFFPOSX1 arr_reg_56__22_ ( .D(n99), .CLK(clk), .Q(arr[1870]) );
  DFFPOSX1 arr_reg_56__21_ ( .D(n85), .CLK(clk), .Q(arr[1869]) );
  DFFPOSX1 arr_reg_56__20_ ( .D(n84), .CLK(clk), .Q(arr[1868]) );
  DFFPOSX1 arr_reg_56__19_ ( .D(n83), .CLK(clk), .Q(arr[1867]) );
  DFFPOSX1 arr_reg_56__18_ ( .D(n82), .CLK(clk), .Q(arr[1866]) );
  DFFPOSX1 arr_reg_56__17_ ( .D(n81), .CLK(clk), .Q(arr[1865]) );
  DFFPOSX1 arr_reg_56__16_ ( .D(n80), .CLK(clk), .Q(arr[1864]) );
  DFFPOSX1 arr_reg_56__15_ ( .D(n79), .CLK(clk), .Q(arr[1863]) );
  DFFPOSX1 arr_reg_56__14_ ( .D(n78), .CLK(clk), .Q(arr[1862]) );
  DFFPOSX1 arr_reg_56__13_ ( .D(n77), .CLK(clk), .Q(arr[1861]) );
  DFFPOSX1 arr_reg_56__12_ ( .D(n76), .CLK(clk), .Q(arr[1860]) );
  DFFPOSX1 arr_reg_56__11_ ( .D(n75), .CLK(clk), .Q(arr[1859]) );
  DFFPOSX1 arr_reg_56__10_ ( .D(n74), .CLK(clk), .Q(arr[1858]) );
  DFFPOSX1 arr_reg_56__9_ ( .D(n73), .CLK(clk), .Q(arr[1857]) );
  DFFPOSX1 arr_reg_56__8_ ( .D(n226), .CLK(clk), .Q(arr[1856]) );
  DFFPOSX1 arr_reg_56__7_ ( .D(n225), .CLK(clk), .Q(arr[1855]) );
  DFFPOSX1 arr_reg_56__6_ ( .D(n72), .CLK(clk), .Q(arr[1854]) );
  DFFPOSX1 arr_reg_56__5_ ( .D(n71), .CLK(clk), .Q(arr[1853]) );
  DFFPOSX1 arr_reg_56__4_ ( .D(n224), .CLK(clk), .Q(arr[1852]) );
  DFFPOSX1 arr_reg_56__3_ ( .D(n223), .CLK(clk), .Q(arr[1851]) );
  DFFPOSX1 arr_reg_56__2_ ( .D(n222), .CLK(clk), .Q(arr[1850]) );
  DFFPOSX1 arr_reg_56__1_ ( .D(n221), .CLK(clk), .Q(arr[1849]) );
  DFFPOSX1 arr_reg_56__0_ ( .D(n220), .CLK(clk), .Q(arr[1848]) );
  DFFPOSX1 arr_reg_55__32_ ( .D(n8605), .CLK(clk), .Q(arr[1847]) );
  DFFPOSX1 arr_reg_55__31_ ( .D(n8604), .CLK(clk), .Q(arr[1846]) );
  DFFPOSX1 arr_reg_55__30_ ( .D(n8603), .CLK(clk), .Q(arr[1845]) );
  DFFPOSX1 arr_reg_55__29_ ( .D(n8602), .CLK(clk), .Q(arr[1844]) );
  DFFPOSX1 arr_reg_55__28_ ( .D(n8601), .CLK(clk), .Q(arr[1843]) );
  DFFPOSX1 arr_reg_55__27_ ( .D(n8600), .CLK(clk), .Q(arr[1842]) );
  DFFPOSX1 arr_reg_55__26_ ( .D(n8599), .CLK(clk), .Q(arr[1841]) );
  DFFPOSX1 arr_reg_55__25_ ( .D(n8598), .CLK(clk), .Q(arr[1840]) );
  DFFPOSX1 arr_reg_55__24_ ( .D(n8597), .CLK(clk), .Q(arr[1839]) );
  DFFPOSX1 arr_reg_55__23_ ( .D(n8596), .CLK(clk), .Q(arr[1838]) );
  DFFPOSX1 arr_reg_55__22_ ( .D(n8595), .CLK(clk), .Q(arr[1837]) );
  DFFPOSX1 arr_reg_55__21_ ( .D(n8594), .CLK(clk), .Q(arr[1836]) );
  DFFPOSX1 arr_reg_55__20_ ( .D(n8593), .CLK(clk), .Q(arr[1835]) );
  DFFPOSX1 arr_reg_55__19_ ( .D(n8592), .CLK(clk), .Q(arr[1834]) );
  DFFPOSX1 arr_reg_55__18_ ( .D(n8591), .CLK(clk), .Q(arr[1833]) );
  DFFPOSX1 arr_reg_55__17_ ( .D(n8590), .CLK(clk), .Q(arr[1832]) );
  DFFPOSX1 arr_reg_55__16_ ( .D(n8589), .CLK(clk), .Q(arr[1831]) );
  DFFPOSX1 arr_reg_55__15_ ( .D(n8588), .CLK(clk), .Q(arr[1830]) );
  DFFPOSX1 arr_reg_55__14_ ( .D(n8587), .CLK(clk), .Q(arr[1829]) );
  DFFPOSX1 arr_reg_55__13_ ( .D(n8586), .CLK(clk), .Q(arr[1828]) );
  DFFPOSX1 arr_reg_55__12_ ( .D(n8585), .CLK(clk), .Q(arr[1827]) );
  DFFPOSX1 arr_reg_55__11_ ( .D(n8584), .CLK(clk), .Q(arr[1826]) );
  DFFPOSX1 arr_reg_55__10_ ( .D(n8583), .CLK(clk), .Q(arr[1825]) );
  DFFPOSX1 arr_reg_55__9_ ( .D(n8582), .CLK(clk), .Q(arr[1824]) );
  DFFPOSX1 arr_reg_55__8_ ( .D(n8581), .CLK(clk), .Q(arr[1823]) );
  DFFPOSX1 arr_reg_55__7_ ( .D(n8580), .CLK(clk), .Q(arr[1822]) );
  DFFPOSX1 arr_reg_55__6_ ( .D(n8579), .CLK(clk), .Q(arr[1821]) );
  DFFPOSX1 arr_reg_55__5_ ( .D(n8578), .CLK(clk), .Q(arr[1820]) );
  DFFPOSX1 arr_reg_55__4_ ( .D(n8577), .CLK(clk), .Q(arr[1819]) );
  DFFPOSX1 arr_reg_55__3_ ( .D(n8576), .CLK(clk), .Q(arr[1818]) );
  DFFPOSX1 arr_reg_55__2_ ( .D(n8575), .CLK(clk), .Q(arr[1817]) );
  DFFPOSX1 arr_reg_55__1_ ( .D(n8574), .CLK(clk), .Q(arr[1816]) );
  DFFPOSX1 arr_reg_55__0_ ( .D(n8573), .CLK(clk), .Q(arr[1815]) );
  DFFPOSX1 arr_reg_54__32_ ( .D(n8572), .CLK(clk), .Q(arr[1814]) );
  DFFPOSX1 arr_reg_54__31_ ( .D(n8571), .CLK(clk), .Q(arr[1813]) );
  DFFPOSX1 arr_reg_54__30_ ( .D(n8570), .CLK(clk), .Q(arr[1812]) );
  DFFPOSX1 arr_reg_54__29_ ( .D(n8569), .CLK(clk), .Q(arr[1811]) );
  DFFPOSX1 arr_reg_54__28_ ( .D(n8568), .CLK(clk), .Q(arr[1810]) );
  DFFPOSX1 arr_reg_54__27_ ( .D(n8567), .CLK(clk), .Q(arr[1809]) );
  DFFPOSX1 arr_reg_54__26_ ( .D(n8566), .CLK(clk), .Q(arr[1808]) );
  DFFPOSX1 arr_reg_54__25_ ( .D(n8565), .CLK(clk), .Q(arr[1807]) );
  DFFPOSX1 arr_reg_54__24_ ( .D(n8564), .CLK(clk), .Q(arr[1806]) );
  DFFPOSX1 arr_reg_54__23_ ( .D(n8563), .CLK(clk), .Q(arr[1805]) );
  DFFPOSX1 arr_reg_54__22_ ( .D(n8562), .CLK(clk), .Q(arr[1804]) );
  DFFPOSX1 arr_reg_54__21_ ( .D(n8561), .CLK(clk), .Q(arr[1803]) );
  DFFPOSX1 arr_reg_54__20_ ( .D(n8560), .CLK(clk), .Q(arr[1802]) );
  DFFPOSX1 arr_reg_54__19_ ( .D(n8559), .CLK(clk), .Q(arr[1801]) );
  DFFPOSX1 arr_reg_54__18_ ( .D(n8558), .CLK(clk), .Q(arr[1800]) );
  DFFPOSX1 arr_reg_54__17_ ( .D(n8557), .CLK(clk), .Q(arr[1799]) );
  DFFPOSX1 arr_reg_54__16_ ( .D(n8556), .CLK(clk), .Q(arr[1798]) );
  DFFPOSX1 arr_reg_54__15_ ( .D(n8555), .CLK(clk), .Q(arr[1797]) );
  DFFPOSX1 arr_reg_54__14_ ( .D(n8554), .CLK(clk), .Q(arr[1796]) );
  DFFPOSX1 arr_reg_54__13_ ( .D(n8553), .CLK(clk), .Q(arr[1795]) );
  DFFPOSX1 arr_reg_54__12_ ( .D(n8552), .CLK(clk), .Q(arr[1794]) );
  DFFPOSX1 arr_reg_54__11_ ( .D(n8551), .CLK(clk), .Q(arr[1793]) );
  DFFPOSX1 arr_reg_54__10_ ( .D(n8550), .CLK(clk), .Q(arr[1792]) );
  DFFPOSX1 arr_reg_54__9_ ( .D(n8549), .CLK(clk), .Q(arr[1791]) );
  DFFPOSX1 arr_reg_54__8_ ( .D(n8548), .CLK(clk), .Q(arr[1790]) );
  DFFPOSX1 arr_reg_54__7_ ( .D(n8547), .CLK(clk), .Q(arr[1789]) );
  DFFPOSX1 arr_reg_54__6_ ( .D(n8546), .CLK(clk), .Q(arr[1788]) );
  DFFPOSX1 arr_reg_54__5_ ( .D(n8545), .CLK(clk), .Q(arr[1787]) );
  DFFPOSX1 arr_reg_54__4_ ( .D(n8544), .CLK(clk), .Q(arr[1786]) );
  DFFPOSX1 arr_reg_54__3_ ( .D(n8543), .CLK(clk), .Q(arr[1785]) );
  DFFPOSX1 arr_reg_54__2_ ( .D(n8542), .CLK(clk), .Q(arr[1784]) );
  DFFPOSX1 arr_reg_54__1_ ( .D(n8541), .CLK(clk), .Q(arr[1783]) );
  DFFPOSX1 arr_reg_54__0_ ( .D(n8540), .CLK(clk), .Q(arr[1782]) );
  DFFPOSX1 arr_reg_53__32_ ( .D(n8539), .CLK(clk), .Q(arr[1781]) );
  DFFPOSX1 arr_reg_53__31_ ( .D(n8538), .CLK(clk), .Q(arr[1780]) );
  DFFPOSX1 arr_reg_53__30_ ( .D(n8537), .CLK(clk), .Q(arr[1779]) );
  DFFPOSX1 arr_reg_53__29_ ( .D(n8536), .CLK(clk), .Q(arr[1778]) );
  DFFPOSX1 arr_reg_53__28_ ( .D(n8535), .CLK(clk), .Q(arr[1777]) );
  DFFPOSX1 arr_reg_53__27_ ( .D(n8534), .CLK(clk), .Q(arr[1776]) );
  DFFPOSX1 arr_reg_53__26_ ( .D(n8533), .CLK(clk), .Q(arr[1775]) );
  DFFPOSX1 arr_reg_53__25_ ( .D(n8532), .CLK(clk), .Q(arr[1774]) );
  DFFPOSX1 arr_reg_53__24_ ( .D(n8531), .CLK(clk), .Q(arr[1773]) );
  DFFPOSX1 arr_reg_53__23_ ( .D(n8530), .CLK(clk), .Q(arr[1772]) );
  DFFPOSX1 arr_reg_53__22_ ( .D(n8529), .CLK(clk), .Q(arr[1771]) );
  DFFPOSX1 arr_reg_53__21_ ( .D(n8528), .CLK(clk), .Q(arr[1770]) );
  DFFPOSX1 arr_reg_53__20_ ( .D(n8527), .CLK(clk), .Q(arr[1769]) );
  DFFPOSX1 arr_reg_53__19_ ( .D(n8526), .CLK(clk), .Q(arr[1768]) );
  DFFPOSX1 arr_reg_53__18_ ( .D(n8525), .CLK(clk), .Q(arr[1767]) );
  DFFPOSX1 arr_reg_53__17_ ( .D(n8524), .CLK(clk), .Q(arr[1766]) );
  DFFPOSX1 arr_reg_53__16_ ( .D(n8523), .CLK(clk), .Q(arr[1765]) );
  DFFPOSX1 arr_reg_53__15_ ( .D(n8522), .CLK(clk), .Q(arr[1764]) );
  DFFPOSX1 arr_reg_53__14_ ( .D(n8521), .CLK(clk), .Q(arr[1763]) );
  DFFPOSX1 arr_reg_53__13_ ( .D(n8520), .CLK(clk), .Q(arr[1762]) );
  DFFPOSX1 arr_reg_53__12_ ( .D(n8519), .CLK(clk), .Q(arr[1761]) );
  DFFPOSX1 arr_reg_53__11_ ( .D(n8518), .CLK(clk), .Q(arr[1760]) );
  DFFPOSX1 arr_reg_53__10_ ( .D(n8517), .CLK(clk), .Q(arr[1759]) );
  DFFPOSX1 arr_reg_53__9_ ( .D(n8516), .CLK(clk), .Q(arr[1758]) );
  DFFPOSX1 arr_reg_53__8_ ( .D(n8515), .CLK(clk), .Q(arr[1757]) );
  DFFPOSX1 arr_reg_53__7_ ( .D(n8514), .CLK(clk), .Q(arr[1756]) );
  DFFPOSX1 arr_reg_53__6_ ( .D(n8513), .CLK(clk), .Q(arr[1755]) );
  DFFPOSX1 arr_reg_53__5_ ( .D(n8512), .CLK(clk), .Q(arr[1754]) );
  DFFPOSX1 arr_reg_53__4_ ( .D(n8511), .CLK(clk), .Q(arr[1753]) );
  DFFPOSX1 arr_reg_53__3_ ( .D(n8510), .CLK(clk), .Q(arr[1752]) );
  DFFPOSX1 arr_reg_53__2_ ( .D(n8509), .CLK(clk), .Q(arr[1751]) );
  DFFPOSX1 arr_reg_53__1_ ( .D(n8508), .CLK(clk), .Q(arr[1750]) );
  DFFPOSX1 arr_reg_53__0_ ( .D(n8507), .CLK(clk), .Q(arr[1749]) );
  DFFPOSX1 arr_reg_52__32_ ( .D(n8506), .CLK(clk), .Q(arr[1748]) );
  DFFPOSX1 arr_reg_52__31_ ( .D(n8505), .CLK(clk), .Q(arr[1747]) );
  DFFPOSX1 arr_reg_52__30_ ( .D(n8504), .CLK(clk), .Q(arr[1746]) );
  DFFPOSX1 arr_reg_52__29_ ( .D(n8503), .CLK(clk), .Q(arr[1745]) );
  DFFPOSX1 arr_reg_52__28_ ( .D(n8502), .CLK(clk), .Q(arr[1744]) );
  DFFPOSX1 arr_reg_52__27_ ( .D(n8501), .CLK(clk), .Q(arr[1743]) );
  DFFPOSX1 arr_reg_52__26_ ( .D(n8500), .CLK(clk), .Q(arr[1742]) );
  DFFPOSX1 arr_reg_52__25_ ( .D(n8499), .CLK(clk), .Q(arr[1741]) );
  DFFPOSX1 arr_reg_52__24_ ( .D(n8498), .CLK(clk), .Q(arr[1740]) );
  DFFPOSX1 arr_reg_52__23_ ( .D(n8497), .CLK(clk), .Q(arr[1739]) );
  DFFPOSX1 arr_reg_52__22_ ( .D(n8496), .CLK(clk), .Q(arr[1738]) );
  DFFPOSX1 arr_reg_52__21_ ( .D(n8495), .CLK(clk), .Q(arr[1737]) );
  DFFPOSX1 arr_reg_52__20_ ( .D(n8494), .CLK(clk), .Q(arr[1736]) );
  DFFPOSX1 arr_reg_52__19_ ( .D(n8493), .CLK(clk), .Q(arr[1735]) );
  DFFPOSX1 arr_reg_52__18_ ( .D(n8492), .CLK(clk), .Q(arr[1734]) );
  DFFPOSX1 arr_reg_52__17_ ( .D(n8491), .CLK(clk), .Q(arr[1733]) );
  DFFPOSX1 arr_reg_52__16_ ( .D(n8490), .CLK(clk), .Q(arr[1732]) );
  DFFPOSX1 arr_reg_52__15_ ( .D(n8489), .CLK(clk), .Q(arr[1731]) );
  DFFPOSX1 arr_reg_52__14_ ( .D(n8488), .CLK(clk), .Q(arr[1730]) );
  DFFPOSX1 arr_reg_52__13_ ( .D(n8487), .CLK(clk), .Q(arr[1729]) );
  DFFPOSX1 arr_reg_52__12_ ( .D(n8486), .CLK(clk), .Q(arr[1728]) );
  DFFPOSX1 arr_reg_52__11_ ( .D(n8485), .CLK(clk), .Q(arr[1727]) );
  DFFPOSX1 arr_reg_52__10_ ( .D(n8484), .CLK(clk), .Q(arr[1726]) );
  DFFPOSX1 arr_reg_52__9_ ( .D(n8483), .CLK(clk), .Q(arr[1725]) );
  DFFPOSX1 arr_reg_52__8_ ( .D(n8482), .CLK(clk), .Q(arr[1724]) );
  DFFPOSX1 arr_reg_52__7_ ( .D(n8481), .CLK(clk), .Q(arr[1723]) );
  DFFPOSX1 arr_reg_52__6_ ( .D(n8480), .CLK(clk), .Q(arr[1722]) );
  DFFPOSX1 arr_reg_52__5_ ( .D(n8479), .CLK(clk), .Q(arr[1721]) );
  DFFPOSX1 arr_reg_52__4_ ( .D(n8478), .CLK(clk), .Q(arr[1720]) );
  DFFPOSX1 arr_reg_52__3_ ( .D(n8477), .CLK(clk), .Q(arr[1719]) );
  DFFPOSX1 arr_reg_52__2_ ( .D(n8476), .CLK(clk), .Q(arr[1718]) );
  DFFPOSX1 arr_reg_52__1_ ( .D(n8475), .CLK(clk), .Q(arr[1717]) );
  DFFPOSX1 arr_reg_52__0_ ( .D(n8474), .CLK(clk), .Q(arr[1716]) );
  DFFPOSX1 arr_reg_51__32_ ( .D(n8473), .CLK(clk), .Q(arr[1715]) );
  DFFPOSX1 arr_reg_51__31_ ( .D(n8472), .CLK(clk), .Q(arr[1714]) );
  DFFPOSX1 arr_reg_51__30_ ( .D(n8471), .CLK(clk), .Q(arr[1713]) );
  DFFPOSX1 arr_reg_51__29_ ( .D(n8470), .CLK(clk), .Q(arr[1712]) );
  DFFPOSX1 arr_reg_51__28_ ( .D(n8469), .CLK(clk), .Q(arr[1711]) );
  DFFPOSX1 arr_reg_51__27_ ( .D(n8468), .CLK(clk), .Q(arr[1710]) );
  DFFPOSX1 arr_reg_51__26_ ( .D(n8467), .CLK(clk), .Q(arr[1709]) );
  DFFPOSX1 arr_reg_51__25_ ( .D(n8466), .CLK(clk), .Q(arr[1708]) );
  DFFPOSX1 arr_reg_51__24_ ( .D(n8465), .CLK(clk), .Q(arr[1707]) );
  DFFPOSX1 arr_reg_51__23_ ( .D(n8464), .CLK(clk), .Q(arr[1706]) );
  DFFPOSX1 arr_reg_51__22_ ( .D(n8463), .CLK(clk), .Q(arr[1705]) );
  DFFPOSX1 arr_reg_51__21_ ( .D(n8462), .CLK(clk), .Q(arr[1704]) );
  DFFPOSX1 arr_reg_51__20_ ( .D(n8461), .CLK(clk), .Q(arr[1703]) );
  DFFPOSX1 arr_reg_51__19_ ( .D(n8460), .CLK(clk), .Q(arr[1702]) );
  DFFPOSX1 arr_reg_51__18_ ( .D(n8459), .CLK(clk), .Q(arr[1701]) );
  DFFPOSX1 arr_reg_51__17_ ( .D(n8458), .CLK(clk), .Q(arr[1700]) );
  DFFPOSX1 arr_reg_51__16_ ( .D(n8457), .CLK(clk), .Q(arr[1699]) );
  DFFPOSX1 arr_reg_51__15_ ( .D(n8456), .CLK(clk), .Q(arr[1698]) );
  DFFPOSX1 arr_reg_51__14_ ( .D(n8455), .CLK(clk), .Q(arr[1697]) );
  DFFPOSX1 arr_reg_51__13_ ( .D(n8454), .CLK(clk), .Q(arr[1696]) );
  DFFPOSX1 arr_reg_51__12_ ( .D(n8453), .CLK(clk), .Q(arr[1695]) );
  DFFPOSX1 arr_reg_51__11_ ( .D(n8452), .CLK(clk), .Q(arr[1694]) );
  DFFPOSX1 arr_reg_51__10_ ( .D(n8451), .CLK(clk), .Q(arr[1693]) );
  DFFPOSX1 arr_reg_51__9_ ( .D(n8450), .CLK(clk), .Q(arr[1692]) );
  DFFPOSX1 arr_reg_51__8_ ( .D(n8449), .CLK(clk), .Q(arr[1691]) );
  DFFPOSX1 arr_reg_51__7_ ( .D(n8448), .CLK(clk), .Q(arr[1690]) );
  DFFPOSX1 arr_reg_51__6_ ( .D(n8447), .CLK(clk), .Q(arr[1689]) );
  DFFPOSX1 arr_reg_51__5_ ( .D(n8446), .CLK(clk), .Q(arr[1688]) );
  DFFPOSX1 arr_reg_51__4_ ( .D(n8445), .CLK(clk), .Q(arr[1687]) );
  DFFPOSX1 arr_reg_51__3_ ( .D(n8444), .CLK(clk), .Q(arr[1686]) );
  DFFPOSX1 arr_reg_51__2_ ( .D(n8443), .CLK(clk), .Q(arr[1685]) );
  DFFPOSX1 arr_reg_51__1_ ( .D(n8442), .CLK(clk), .Q(arr[1684]) );
  DFFPOSX1 arr_reg_51__0_ ( .D(n8441), .CLK(clk), .Q(arr[1683]) );
  DFFPOSX1 arr_reg_50__32_ ( .D(n8440), .CLK(clk), .Q(arr[1682]) );
  DFFPOSX1 arr_reg_50__31_ ( .D(n8439), .CLK(clk), .Q(arr[1681]) );
  DFFPOSX1 arr_reg_50__30_ ( .D(n8438), .CLK(clk), .Q(arr[1680]) );
  DFFPOSX1 arr_reg_50__29_ ( .D(n8437), .CLK(clk), .Q(arr[1679]) );
  DFFPOSX1 arr_reg_50__28_ ( .D(n8436), .CLK(clk), .Q(arr[1678]) );
  DFFPOSX1 arr_reg_50__27_ ( .D(n8435), .CLK(clk), .Q(arr[1677]) );
  DFFPOSX1 arr_reg_50__26_ ( .D(n8434), .CLK(clk), .Q(arr[1676]) );
  DFFPOSX1 arr_reg_50__25_ ( .D(n8433), .CLK(clk), .Q(arr[1675]) );
  DFFPOSX1 arr_reg_50__24_ ( .D(n8432), .CLK(clk), .Q(arr[1674]) );
  DFFPOSX1 arr_reg_50__23_ ( .D(n8431), .CLK(clk), .Q(arr[1673]) );
  DFFPOSX1 arr_reg_50__22_ ( .D(n8430), .CLK(clk), .Q(arr[1672]) );
  DFFPOSX1 arr_reg_50__21_ ( .D(n8429), .CLK(clk), .Q(arr[1671]) );
  DFFPOSX1 arr_reg_50__20_ ( .D(n8428), .CLK(clk), .Q(arr[1670]) );
  DFFPOSX1 arr_reg_50__19_ ( .D(n8427), .CLK(clk), .Q(arr[1669]) );
  DFFPOSX1 arr_reg_50__18_ ( .D(n8426), .CLK(clk), .Q(arr[1668]) );
  DFFPOSX1 arr_reg_50__17_ ( .D(n8425), .CLK(clk), .Q(arr[1667]) );
  DFFPOSX1 arr_reg_50__16_ ( .D(n8424), .CLK(clk), .Q(arr[1666]) );
  DFFPOSX1 arr_reg_50__15_ ( .D(n8423), .CLK(clk), .Q(arr[1665]) );
  DFFPOSX1 arr_reg_50__14_ ( .D(n8422), .CLK(clk), .Q(arr[1664]) );
  DFFPOSX1 arr_reg_50__13_ ( .D(n8421), .CLK(clk), .Q(arr[1663]) );
  DFFPOSX1 arr_reg_50__12_ ( .D(n8420), .CLK(clk), .Q(arr[1662]) );
  DFFPOSX1 arr_reg_50__11_ ( .D(n8419), .CLK(clk), .Q(arr[1661]) );
  DFFPOSX1 arr_reg_50__10_ ( .D(n8418), .CLK(clk), .Q(arr[1660]) );
  DFFPOSX1 arr_reg_50__9_ ( .D(n8417), .CLK(clk), .Q(arr[1659]) );
  DFFPOSX1 arr_reg_50__8_ ( .D(n8416), .CLK(clk), .Q(arr[1658]) );
  DFFPOSX1 arr_reg_50__7_ ( .D(n8415), .CLK(clk), .Q(arr[1657]) );
  DFFPOSX1 arr_reg_50__6_ ( .D(n8414), .CLK(clk), .Q(arr[1656]) );
  DFFPOSX1 arr_reg_50__5_ ( .D(n8413), .CLK(clk), .Q(arr[1655]) );
  DFFPOSX1 arr_reg_50__4_ ( .D(n8412), .CLK(clk), .Q(arr[1654]) );
  DFFPOSX1 arr_reg_50__3_ ( .D(n8411), .CLK(clk), .Q(arr[1653]) );
  DFFPOSX1 arr_reg_50__2_ ( .D(n8410), .CLK(clk), .Q(arr[1652]) );
  DFFPOSX1 arr_reg_50__1_ ( .D(n8409), .CLK(clk), .Q(arr[1651]) );
  DFFPOSX1 arr_reg_50__0_ ( .D(n8408), .CLK(clk), .Q(arr[1650]) );
  DFFPOSX1 arr_reg_49__32_ ( .D(n8407), .CLK(clk), .Q(arr[1649]) );
  DFFPOSX1 arr_reg_49__31_ ( .D(n8406), .CLK(clk), .Q(arr[1648]) );
  DFFPOSX1 arr_reg_49__30_ ( .D(n8405), .CLK(clk), .Q(arr[1647]) );
  DFFPOSX1 arr_reg_49__29_ ( .D(n8404), .CLK(clk), .Q(arr[1646]) );
  DFFPOSX1 arr_reg_49__28_ ( .D(n8403), .CLK(clk), .Q(arr[1645]) );
  DFFPOSX1 arr_reg_49__27_ ( .D(n8402), .CLK(clk), .Q(arr[1644]) );
  DFFPOSX1 arr_reg_49__26_ ( .D(n8401), .CLK(clk), .Q(arr[1643]) );
  DFFPOSX1 arr_reg_49__25_ ( .D(n8400), .CLK(clk), .Q(arr[1642]) );
  DFFPOSX1 arr_reg_49__24_ ( .D(n8399), .CLK(clk), .Q(arr[1641]) );
  DFFPOSX1 arr_reg_49__23_ ( .D(n8398), .CLK(clk), .Q(arr[1640]) );
  DFFPOSX1 arr_reg_49__22_ ( .D(n8397), .CLK(clk), .Q(arr[1639]) );
  DFFPOSX1 arr_reg_49__21_ ( .D(n8396), .CLK(clk), .Q(arr[1638]) );
  DFFPOSX1 arr_reg_49__20_ ( .D(n8395), .CLK(clk), .Q(arr[1637]) );
  DFFPOSX1 arr_reg_49__19_ ( .D(n8394), .CLK(clk), .Q(arr[1636]) );
  DFFPOSX1 arr_reg_49__18_ ( .D(n8393), .CLK(clk), .Q(arr[1635]) );
  DFFPOSX1 arr_reg_49__17_ ( .D(n8392), .CLK(clk), .Q(arr[1634]) );
  DFFPOSX1 arr_reg_49__16_ ( .D(n8391), .CLK(clk), .Q(arr[1633]) );
  DFFPOSX1 arr_reg_49__15_ ( .D(n8390), .CLK(clk), .Q(arr[1632]) );
  DFFPOSX1 arr_reg_49__14_ ( .D(n8389), .CLK(clk), .Q(arr[1631]) );
  DFFPOSX1 arr_reg_49__13_ ( .D(n8388), .CLK(clk), .Q(arr[1630]) );
  DFFPOSX1 arr_reg_49__12_ ( .D(n8387), .CLK(clk), .Q(arr[1629]) );
  DFFPOSX1 arr_reg_49__11_ ( .D(n8386), .CLK(clk), .Q(arr[1628]) );
  DFFPOSX1 arr_reg_49__10_ ( .D(n8385), .CLK(clk), .Q(arr[1627]) );
  DFFPOSX1 arr_reg_49__9_ ( .D(n8384), .CLK(clk), .Q(arr[1626]) );
  DFFPOSX1 arr_reg_49__8_ ( .D(n8383), .CLK(clk), .Q(arr[1625]) );
  DFFPOSX1 arr_reg_49__7_ ( .D(n8382), .CLK(clk), .Q(arr[1624]) );
  DFFPOSX1 arr_reg_49__6_ ( .D(n8381), .CLK(clk), .Q(arr[1623]) );
  DFFPOSX1 arr_reg_49__5_ ( .D(n8380), .CLK(clk), .Q(arr[1622]) );
  DFFPOSX1 arr_reg_49__4_ ( .D(n8379), .CLK(clk), .Q(arr[1621]) );
  DFFPOSX1 arr_reg_49__3_ ( .D(n8378), .CLK(clk), .Q(arr[1620]) );
  DFFPOSX1 arr_reg_49__2_ ( .D(n8377), .CLK(clk), .Q(arr[1619]) );
  DFFPOSX1 arr_reg_49__1_ ( .D(n8376), .CLK(clk), .Q(arr[1618]) );
  DFFPOSX1 arr_reg_49__0_ ( .D(n8375), .CLK(clk), .Q(arr[1617]) );
  DFFPOSX1 arr_reg_48__32_ ( .D(n8374), .CLK(clk), .Q(arr[1616]) );
  DFFPOSX1 arr_reg_48__31_ ( .D(n8373), .CLK(clk), .Q(arr[1615]) );
  DFFPOSX1 arr_reg_48__30_ ( .D(n8372), .CLK(clk), .Q(arr[1614]) );
  DFFPOSX1 arr_reg_48__29_ ( .D(n8371), .CLK(clk), .Q(arr[1613]) );
  DFFPOSX1 arr_reg_48__28_ ( .D(n8370), .CLK(clk), .Q(arr[1612]) );
  DFFPOSX1 arr_reg_48__27_ ( .D(n8369), .CLK(clk), .Q(arr[1611]) );
  DFFPOSX1 arr_reg_48__26_ ( .D(n8368), .CLK(clk), .Q(arr[1610]) );
  DFFPOSX1 arr_reg_48__25_ ( .D(n8367), .CLK(clk), .Q(arr[1609]) );
  DFFPOSX1 arr_reg_48__24_ ( .D(n8366), .CLK(clk), .Q(arr[1608]) );
  DFFPOSX1 arr_reg_48__23_ ( .D(n8365), .CLK(clk), .Q(arr[1607]) );
  DFFPOSX1 arr_reg_48__22_ ( .D(n8364), .CLK(clk), .Q(arr[1606]) );
  DFFPOSX1 arr_reg_48__21_ ( .D(n8363), .CLK(clk), .Q(arr[1605]) );
  DFFPOSX1 arr_reg_48__20_ ( .D(n8362), .CLK(clk), .Q(arr[1604]) );
  DFFPOSX1 arr_reg_48__19_ ( .D(n8361), .CLK(clk), .Q(arr[1603]) );
  DFFPOSX1 arr_reg_48__18_ ( .D(n8360), .CLK(clk), .Q(arr[1602]) );
  DFFPOSX1 arr_reg_48__17_ ( .D(n8359), .CLK(clk), .Q(arr[1601]) );
  DFFPOSX1 arr_reg_48__16_ ( .D(n8358), .CLK(clk), .Q(arr[1600]) );
  DFFPOSX1 arr_reg_48__15_ ( .D(n8357), .CLK(clk), .Q(arr[1599]) );
  DFFPOSX1 arr_reg_48__14_ ( .D(n8356), .CLK(clk), .Q(arr[1598]) );
  DFFPOSX1 arr_reg_48__13_ ( .D(n8355), .CLK(clk), .Q(arr[1597]) );
  DFFPOSX1 arr_reg_48__12_ ( .D(n8354), .CLK(clk), .Q(arr[1596]) );
  DFFPOSX1 arr_reg_48__11_ ( .D(n8353), .CLK(clk), .Q(arr[1595]) );
  DFFPOSX1 arr_reg_48__10_ ( .D(n8352), .CLK(clk), .Q(arr[1594]) );
  DFFPOSX1 arr_reg_48__9_ ( .D(n8351), .CLK(clk), .Q(arr[1593]) );
  DFFPOSX1 arr_reg_48__8_ ( .D(n8350), .CLK(clk), .Q(arr[1592]) );
  DFFPOSX1 arr_reg_48__7_ ( .D(n8349), .CLK(clk), .Q(arr[1591]) );
  DFFPOSX1 arr_reg_48__6_ ( .D(n8348), .CLK(clk), .Q(arr[1590]) );
  DFFPOSX1 arr_reg_48__5_ ( .D(n8347), .CLK(clk), .Q(arr[1589]) );
  DFFPOSX1 arr_reg_48__4_ ( .D(n8346), .CLK(clk), .Q(arr[1588]) );
  DFFPOSX1 arr_reg_48__3_ ( .D(n8345), .CLK(clk), .Q(arr[1587]) );
  DFFPOSX1 arr_reg_48__2_ ( .D(n8344), .CLK(clk), .Q(arr[1586]) );
  DFFPOSX1 arr_reg_48__1_ ( .D(n8343), .CLK(clk), .Q(arr[1585]) );
  DFFPOSX1 arr_reg_48__0_ ( .D(n8342), .CLK(clk), .Q(arr[1584]) );
  DFFPOSX1 arr_reg_47__32_ ( .D(n8341), .CLK(clk), .Q(arr[1583]) );
  DFFPOSX1 arr_reg_47__31_ ( .D(n8340), .CLK(clk), .Q(arr[1582]) );
  DFFPOSX1 arr_reg_47__30_ ( .D(n8339), .CLK(clk), .Q(arr[1581]) );
  DFFPOSX1 arr_reg_47__29_ ( .D(n8338), .CLK(clk), .Q(arr[1580]) );
  DFFPOSX1 arr_reg_47__28_ ( .D(n8337), .CLK(clk), .Q(arr[1579]) );
  DFFPOSX1 arr_reg_47__27_ ( .D(n8336), .CLK(clk), .Q(arr[1578]) );
  DFFPOSX1 arr_reg_47__26_ ( .D(n8335), .CLK(clk), .Q(arr[1577]) );
  DFFPOSX1 arr_reg_47__25_ ( .D(n8334), .CLK(clk), .Q(arr[1576]) );
  DFFPOSX1 arr_reg_47__24_ ( .D(n8333), .CLK(clk), .Q(arr[1575]) );
  DFFPOSX1 arr_reg_47__23_ ( .D(n8332), .CLK(clk), .Q(arr[1574]) );
  DFFPOSX1 arr_reg_47__22_ ( .D(n8331), .CLK(clk), .Q(arr[1573]) );
  DFFPOSX1 arr_reg_47__21_ ( .D(n8330), .CLK(clk), .Q(arr[1572]) );
  DFFPOSX1 arr_reg_47__20_ ( .D(n8329), .CLK(clk), .Q(arr[1571]) );
  DFFPOSX1 arr_reg_47__19_ ( .D(n8328), .CLK(clk), .Q(arr[1570]) );
  DFFPOSX1 arr_reg_47__18_ ( .D(n8327), .CLK(clk), .Q(arr[1569]) );
  DFFPOSX1 arr_reg_47__17_ ( .D(n8326), .CLK(clk), .Q(arr[1568]) );
  DFFPOSX1 arr_reg_47__16_ ( .D(n8325), .CLK(clk), .Q(arr[1567]) );
  DFFPOSX1 arr_reg_47__15_ ( .D(n8324), .CLK(clk), .Q(arr[1566]) );
  DFFPOSX1 arr_reg_47__14_ ( .D(n8323), .CLK(clk), .Q(arr[1565]) );
  DFFPOSX1 arr_reg_47__13_ ( .D(n8322), .CLK(clk), .Q(arr[1564]) );
  DFFPOSX1 arr_reg_47__12_ ( .D(n8321), .CLK(clk), .Q(arr[1563]) );
  DFFPOSX1 arr_reg_47__11_ ( .D(n8320), .CLK(clk), .Q(arr[1562]) );
  DFFPOSX1 arr_reg_47__10_ ( .D(n8319), .CLK(clk), .Q(arr[1561]) );
  DFFPOSX1 arr_reg_47__9_ ( .D(n8318), .CLK(clk), .Q(arr[1560]) );
  DFFPOSX1 arr_reg_47__8_ ( .D(n8317), .CLK(clk), .Q(arr[1559]) );
  DFFPOSX1 arr_reg_47__7_ ( .D(n8316), .CLK(clk), .Q(arr[1558]) );
  DFFPOSX1 arr_reg_47__6_ ( .D(n8315), .CLK(clk), .Q(arr[1557]) );
  DFFPOSX1 arr_reg_47__5_ ( .D(n8314), .CLK(clk), .Q(arr[1556]) );
  DFFPOSX1 arr_reg_47__4_ ( .D(n8313), .CLK(clk), .Q(arr[1555]) );
  DFFPOSX1 arr_reg_47__3_ ( .D(n8312), .CLK(clk), .Q(arr[1554]) );
  DFFPOSX1 arr_reg_47__2_ ( .D(n8311), .CLK(clk), .Q(arr[1553]) );
  DFFPOSX1 arr_reg_47__1_ ( .D(n8310), .CLK(clk), .Q(arr[1552]) );
  DFFPOSX1 arr_reg_47__0_ ( .D(n8309), .CLK(clk), .Q(arr[1551]) );
  DFFPOSX1 arr_reg_46__32_ ( .D(n8308), .CLK(clk), .Q(arr[1550]) );
  DFFPOSX1 arr_reg_46__31_ ( .D(n8307), .CLK(clk), .Q(arr[1549]) );
  DFFPOSX1 arr_reg_46__30_ ( .D(n8306), .CLK(clk), .Q(arr[1548]) );
  DFFPOSX1 arr_reg_46__29_ ( .D(n8305), .CLK(clk), .Q(arr[1547]) );
  DFFPOSX1 arr_reg_46__28_ ( .D(n8304), .CLK(clk), .Q(arr[1546]) );
  DFFPOSX1 arr_reg_46__27_ ( .D(n8303), .CLK(clk), .Q(arr[1545]) );
  DFFPOSX1 arr_reg_46__26_ ( .D(n8302), .CLK(clk), .Q(arr[1544]) );
  DFFPOSX1 arr_reg_46__25_ ( .D(n8301), .CLK(clk), .Q(arr[1543]) );
  DFFPOSX1 arr_reg_46__24_ ( .D(n8300), .CLK(clk), .Q(arr[1542]) );
  DFFPOSX1 arr_reg_46__23_ ( .D(n8299), .CLK(clk), .Q(arr[1541]) );
  DFFPOSX1 arr_reg_46__22_ ( .D(n8298), .CLK(clk), .Q(arr[1540]) );
  DFFPOSX1 arr_reg_46__21_ ( .D(n8297), .CLK(clk), .Q(arr[1539]) );
  DFFPOSX1 arr_reg_46__20_ ( .D(n8296), .CLK(clk), .Q(arr[1538]) );
  DFFPOSX1 arr_reg_46__19_ ( .D(n8295), .CLK(clk), .Q(arr[1537]) );
  DFFPOSX1 arr_reg_46__18_ ( .D(n8294), .CLK(clk), .Q(arr[1536]) );
  DFFPOSX1 arr_reg_46__17_ ( .D(n8293), .CLK(clk), .Q(arr[1535]) );
  DFFPOSX1 arr_reg_46__16_ ( .D(n8292), .CLK(clk), .Q(arr[1534]) );
  DFFPOSX1 arr_reg_46__15_ ( .D(n8291), .CLK(clk), .Q(arr[1533]) );
  DFFPOSX1 arr_reg_46__14_ ( .D(n8290), .CLK(clk), .Q(arr[1532]) );
  DFFPOSX1 arr_reg_46__13_ ( .D(n8289), .CLK(clk), .Q(arr[1531]) );
  DFFPOSX1 arr_reg_46__12_ ( .D(n8288), .CLK(clk), .Q(arr[1530]) );
  DFFPOSX1 arr_reg_46__11_ ( .D(n8287), .CLK(clk), .Q(arr[1529]) );
  DFFPOSX1 arr_reg_46__10_ ( .D(n8286), .CLK(clk), .Q(arr[1528]) );
  DFFPOSX1 arr_reg_46__9_ ( .D(n8285), .CLK(clk), .Q(arr[1527]) );
  DFFPOSX1 arr_reg_46__8_ ( .D(n8284), .CLK(clk), .Q(arr[1526]) );
  DFFPOSX1 arr_reg_46__7_ ( .D(n8283), .CLK(clk), .Q(arr[1525]) );
  DFFPOSX1 arr_reg_46__6_ ( .D(n8282), .CLK(clk), .Q(arr[1524]) );
  DFFPOSX1 arr_reg_46__5_ ( .D(n8281), .CLK(clk), .Q(arr[1523]) );
  DFFPOSX1 arr_reg_46__4_ ( .D(n8280), .CLK(clk), .Q(arr[1522]) );
  DFFPOSX1 arr_reg_46__3_ ( .D(n8279), .CLK(clk), .Q(arr[1521]) );
  DFFPOSX1 arr_reg_46__2_ ( .D(n8278), .CLK(clk), .Q(arr[1520]) );
  DFFPOSX1 arr_reg_46__1_ ( .D(n8277), .CLK(clk), .Q(arr[1519]) );
  DFFPOSX1 arr_reg_46__0_ ( .D(n8276), .CLK(clk), .Q(arr[1518]) );
  DFFPOSX1 arr_reg_45__32_ ( .D(n8275), .CLK(clk), .Q(arr[1517]) );
  DFFPOSX1 arr_reg_45__31_ ( .D(n8274), .CLK(clk), .Q(arr[1516]) );
  DFFPOSX1 arr_reg_45__30_ ( .D(n8273), .CLK(clk), .Q(arr[1515]) );
  DFFPOSX1 arr_reg_45__29_ ( .D(n8272), .CLK(clk), .Q(arr[1514]) );
  DFFPOSX1 arr_reg_45__28_ ( .D(n8271), .CLK(clk), .Q(arr[1513]) );
  DFFPOSX1 arr_reg_45__27_ ( .D(n8270), .CLK(clk), .Q(arr[1512]) );
  DFFPOSX1 arr_reg_45__26_ ( .D(n8269), .CLK(clk), .Q(arr[1511]) );
  DFFPOSX1 arr_reg_45__25_ ( .D(n8268), .CLK(clk), .Q(arr[1510]) );
  DFFPOSX1 arr_reg_45__24_ ( .D(n8267), .CLK(clk), .Q(arr[1509]) );
  DFFPOSX1 arr_reg_45__23_ ( .D(n8266), .CLK(clk), .Q(arr[1508]) );
  DFFPOSX1 arr_reg_45__22_ ( .D(n8265), .CLK(clk), .Q(arr[1507]) );
  DFFPOSX1 arr_reg_45__21_ ( .D(n8264), .CLK(clk), .Q(arr[1506]) );
  DFFPOSX1 arr_reg_45__20_ ( .D(n8263), .CLK(clk), .Q(arr[1505]) );
  DFFPOSX1 arr_reg_45__19_ ( .D(n8262), .CLK(clk), .Q(arr[1504]) );
  DFFPOSX1 arr_reg_45__18_ ( .D(n8261), .CLK(clk), .Q(arr[1503]) );
  DFFPOSX1 arr_reg_45__17_ ( .D(n8260), .CLK(clk), .Q(arr[1502]) );
  DFFPOSX1 arr_reg_45__16_ ( .D(n8259), .CLK(clk), .Q(arr[1501]) );
  DFFPOSX1 arr_reg_45__15_ ( .D(n8258), .CLK(clk), .Q(arr[1500]) );
  DFFPOSX1 arr_reg_45__14_ ( .D(n8257), .CLK(clk), .Q(arr[1499]) );
  DFFPOSX1 arr_reg_45__13_ ( .D(n8256), .CLK(clk), .Q(arr[1498]) );
  DFFPOSX1 arr_reg_45__12_ ( .D(n8255), .CLK(clk), .Q(arr[1497]) );
  DFFPOSX1 arr_reg_45__11_ ( .D(n8254), .CLK(clk), .Q(arr[1496]) );
  DFFPOSX1 arr_reg_45__10_ ( .D(n8253), .CLK(clk), .Q(arr[1495]) );
  DFFPOSX1 arr_reg_45__9_ ( .D(n8252), .CLK(clk), .Q(arr[1494]) );
  DFFPOSX1 arr_reg_45__8_ ( .D(n8251), .CLK(clk), .Q(arr[1493]) );
  DFFPOSX1 arr_reg_45__7_ ( .D(n8250), .CLK(clk), .Q(arr[1492]) );
  DFFPOSX1 arr_reg_45__6_ ( .D(n8249), .CLK(clk), .Q(arr[1491]) );
  DFFPOSX1 arr_reg_45__5_ ( .D(n8248), .CLK(clk), .Q(arr[1490]) );
  DFFPOSX1 arr_reg_45__4_ ( .D(n8247), .CLK(clk), .Q(arr[1489]) );
  DFFPOSX1 arr_reg_45__3_ ( .D(n8246), .CLK(clk), .Q(arr[1488]) );
  DFFPOSX1 arr_reg_45__2_ ( .D(n8245), .CLK(clk), .Q(arr[1487]) );
  DFFPOSX1 arr_reg_45__1_ ( .D(n8244), .CLK(clk), .Q(arr[1486]) );
  DFFPOSX1 arr_reg_45__0_ ( .D(n8243), .CLK(clk), .Q(arr[1485]) );
  DFFPOSX1 arr_reg_44__32_ ( .D(n8242), .CLK(clk), .Q(arr[1484]) );
  DFFPOSX1 arr_reg_44__31_ ( .D(n8241), .CLK(clk), .Q(arr[1483]) );
  DFFPOSX1 arr_reg_44__30_ ( .D(n8240), .CLK(clk), .Q(arr[1482]) );
  DFFPOSX1 arr_reg_44__29_ ( .D(n8239), .CLK(clk), .Q(arr[1481]) );
  DFFPOSX1 arr_reg_44__28_ ( .D(n8238), .CLK(clk), .Q(arr[1480]) );
  DFFPOSX1 arr_reg_44__27_ ( .D(n8237), .CLK(clk), .Q(arr[1479]) );
  DFFPOSX1 arr_reg_44__26_ ( .D(n8236), .CLK(clk), .Q(arr[1478]) );
  DFFPOSX1 arr_reg_44__25_ ( .D(n8235), .CLK(clk), .Q(arr[1477]) );
  DFFPOSX1 arr_reg_44__24_ ( .D(n8234), .CLK(clk), .Q(arr[1476]) );
  DFFPOSX1 arr_reg_44__23_ ( .D(n8233), .CLK(clk), .Q(arr[1475]) );
  DFFPOSX1 arr_reg_44__22_ ( .D(n8232), .CLK(clk), .Q(arr[1474]) );
  DFFPOSX1 arr_reg_44__21_ ( .D(n8231), .CLK(clk), .Q(arr[1473]) );
  DFFPOSX1 arr_reg_44__20_ ( .D(n8230), .CLK(clk), .Q(arr[1472]) );
  DFFPOSX1 arr_reg_44__19_ ( .D(n8229), .CLK(clk), .Q(arr[1471]) );
  DFFPOSX1 arr_reg_44__18_ ( .D(n8228), .CLK(clk), .Q(arr[1470]) );
  DFFPOSX1 arr_reg_44__17_ ( .D(n8227), .CLK(clk), .Q(arr[1469]) );
  DFFPOSX1 arr_reg_44__16_ ( .D(n8226), .CLK(clk), .Q(arr[1468]) );
  DFFPOSX1 arr_reg_44__15_ ( .D(n8225), .CLK(clk), .Q(arr[1467]) );
  DFFPOSX1 arr_reg_44__14_ ( .D(n8224), .CLK(clk), .Q(arr[1466]) );
  DFFPOSX1 arr_reg_44__13_ ( .D(n8223), .CLK(clk), .Q(arr[1465]) );
  DFFPOSX1 arr_reg_44__12_ ( .D(n8222), .CLK(clk), .Q(arr[1464]) );
  DFFPOSX1 arr_reg_44__11_ ( .D(n8221), .CLK(clk), .Q(arr[1463]) );
  DFFPOSX1 arr_reg_44__10_ ( .D(n8220), .CLK(clk), .Q(arr[1462]) );
  DFFPOSX1 arr_reg_44__9_ ( .D(n8219), .CLK(clk), .Q(arr[1461]) );
  DFFPOSX1 arr_reg_44__8_ ( .D(n8218), .CLK(clk), .Q(arr[1460]) );
  DFFPOSX1 arr_reg_44__7_ ( .D(n8217), .CLK(clk), .Q(arr[1459]) );
  DFFPOSX1 arr_reg_44__6_ ( .D(n8216), .CLK(clk), .Q(arr[1458]) );
  DFFPOSX1 arr_reg_44__5_ ( .D(n8215), .CLK(clk), .Q(arr[1457]) );
  DFFPOSX1 arr_reg_44__4_ ( .D(n8214), .CLK(clk), .Q(arr[1456]) );
  DFFPOSX1 arr_reg_44__3_ ( .D(n8213), .CLK(clk), .Q(arr[1455]) );
  DFFPOSX1 arr_reg_44__2_ ( .D(n8212), .CLK(clk), .Q(arr[1454]) );
  DFFPOSX1 arr_reg_44__1_ ( .D(n8211), .CLK(clk), .Q(arr[1453]) );
  DFFPOSX1 arr_reg_44__0_ ( .D(n8210), .CLK(clk), .Q(arr[1452]) );
  DFFPOSX1 arr_reg_43__32_ ( .D(n8209), .CLK(clk), .Q(arr[1451]) );
  DFFPOSX1 arr_reg_43__31_ ( .D(n8208), .CLK(clk), .Q(arr[1450]) );
  DFFPOSX1 arr_reg_43__30_ ( .D(n8207), .CLK(clk), .Q(arr[1449]) );
  DFFPOSX1 arr_reg_43__29_ ( .D(n8206), .CLK(clk), .Q(arr[1448]) );
  DFFPOSX1 arr_reg_43__28_ ( .D(n8205), .CLK(clk), .Q(arr[1447]) );
  DFFPOSX1 arr_reg_43__27_ ( .D(n8204), .CLK(clk), .Q(arr[1446]) );
  DFFPOSX1 arr_reg_43__26_ ( .D(n8203), .CLK(clk), .Q(arr[1445]) );
  DFFPOSX1 arr_reg_43__25_ ( .D(n8202), .CLK(clk), .Q(arr[1444]) );
  DFFPOSX1 arr_reg_43__24_ ( .D(n8201), .CLK(clk), .Q(arr[1443]) );
  DFFPOSX1 arr_reg_43__23_ ( .D(n8200), .CLK(clk), .Q(arr[1442]) );
  DFFPOSX1 arr_reg_43__22_ ( .D(n8199), .CLK(clk), .Q(arr[1441]) );
  DFFPOSX1 arr_reg_43__21_ ( .D(n8198), .CLK(clk), .Q(arr[1440]) );
  DFFPOSX1 arr_reg_43__20_ ( .D(n8197), .CLK(clk), .Q(arr[1439]) );
  DFFPOSX1 arr_reg_43__19_ ( .D(n8196), .CLK(clk), .Q(arr[1438]) );
  DFFPOSX1 arr_reg_43__18_ ( .D(n8195), .CLK(clk), .Q(arr[1437]) );
  DFFPOSX1 arr_reg_43__17_ ( .D(n8194), .CLK(clk), .Q(arr[1436]) );
  DFFPOSX1 arr_reg_43__16_ ( .D(n8193), .CLK(clk), .Q(arr[1435]) );
  DFFPOSX1 arr_reg_43__15_ ( .D(n8192), .CLK(clk), .Q(arr[1434]) );
  DFFPOSX1 arr_reg_43__14_ ( .D(n8191), .CLK(clk), .Q(arr[1433]) );
  DFFPOSX1 arr_reg_43__13_ ( .D(n8190), .CLK(clk), .Q(arr[1432]) );
  DFFPOSX1 arr_reg_43__12_ ( .D(n8189), .CLK(clk), .Q(arr[1431]) );
  DFFPOSX1 arr_reg_43__11_ ( .D(n8188), .CLK(clk), .Q(arr[1430]) );
  DFFPOSX1 arr_reg_43__10_ ( .D(n8187), .CLK(clk), .Q(arr[1429]) );
  DFFPOSX1 arr_reg_43__9_ ( .D(n8186), .CLK(clk), .Q(arr[1428]) );
  DFFPOSX1 arr_reg_43__8_ ( .D(n8185), .CLK(clk), .Q(arr[1427]) );
  DFFPOSX1 arr_reg_43__7_ ( .D(n8184), .CLK(clk), .Q(arr[1426]) );
  DFFPOSX1 arr_reg_43__6_ ( .D(n8183), .CLK(clk), .Q(arr[1425]) );
  DFFPOSX1 arr_reg_43__5_ ( .D(n8182), .CLK(clk), .Q(arr[1424]) );
  DFFPOSX1 arr_reg_43__4_ ( .D(n8181), .CLK(clk), .Q(arr[1423]) );
  DFFPOSX1 arr_reg_43__3_ ( .D(n8180), .CLK(clk), .Q(arr[1422]) );
  DFFPOSX1 arr_reg_43__2_ ( .D(n8179), .CLK(clk), .Q(arr[1421]) );
  DFFPOSX1 arr_reg_43__1_ ( .D(n8178), .CLK(clk), .Q(arr[1420]) );
  DFFPOSX1 arr_reg_43__0_ ( .D(n8177), .CLK(clk), .Q(arr[1419]) );
  DFFPOSX1 arr_reg_42__32_ ( .D(n8176), .CLK(clk), .Q(arr[1418]) );
  DFFPOSX1 arr_reg_42__31_ ( .D(n8175), .CLK(clk), .Q(arr[1417]) );
  DFFPOSX1 arr_reg_42__30_ ( .D(n8174), .CLK(clk), .Q(arr[1416]) );
  DFFPOSX1 arr_reg_42__29_ ( .D(n8173), .CLK(clk), .Q(arr[1415]) );
  DFFPOSX1 arr_reg_42__28_ ( .D(n8172), .CLK(clk), .Q(arr[1414]) );
  DFFPOSX1 arr_reg_42__27_ ( .D(n8171), .CLK(clk), .Q(arr[1413]) );
  DFFPOSX1 arr_reg_42__26_ ( .D(n8170), .CLK(clk), .Q(arr[1412]) );
  DFFPOSX1 arr_reg_42__25_ ( .D(n8169), .CLK(clk), .Q(arr[1411]) );
  DFFPOSX1 arr_reg_42__24_ ( .D(n8168), .CLK(clk), .Q(arr[1410]) );
  DFFPOSX1 arr_reg_42__23_ ( .D(n8167), .CLK(clk), .Q(arr[1409]) );
  DFFPOSX1 arr_reg_42__22_ ( .D(n8166), .CLK(clk), .Q(arr[1408]) );
  DFFPOSX1 arr_reg_42__21_ ( .D(n8165), .CLK(clk), .Q(arr[1407]) );
  DFFPOSX1 arr_reg_42__20_ ( .D(n8164), .CLK(clk), .Q(arr[1406]) );
  DFFPOSX1 arr_reg_42__19_ ( .D(n8163), .CLK(clk), .Q(arr[1405]) );
  DFFPOSX1 arr_reg_42__18_ ( .D(n8162), .CLK(clk), .Q(arr[1404]) );
  DFFPOSX1 arr_reg_42__17_ ( .D(n8161), .CLK(clk), .Q(arr[1403]) );
  DFFPOSX1 arr_reg_42__16_ ( .D(n8160), .CLK(clk), .Q(arr[1402]) );
  DFFPOSX1 arr_reg_42__15_ ( .D(n8159), .CLK(clk), .Q(arr[1401]) );
  DFFPOSX1 arr_reg_42__14_ ( .D(n8158), .CLK(clk), .Q(arr[1400]) );
  DFFPOSX1 arr_reg_42__13_ ( .D(n8157), .CLK(clk), .Q(arr[1399]) );
  DFFPOSX1 arr_reg_42__12_ ( .D(n8156), .CLK(clk), .Q(arr[1398]) );
  DFFPOSX1 arr_reg_42__11_ ( .D(n8155), .CLK(clk), .Q(arr[1397]) );
  DFFPOSX1 arr_reg_42__10_ ( .D(n8154), .CLK(clk), .Q(arr[1396]) );
  DFFPOSX1 arr_reg_42__9_ ( .D(n8153), .CLK(clk), .Q(arr[1395]) );
  DFFPOSX1 arr_reg_42__8_ ( .D(n8152), .CLK(clk), .Q(arr[1394]) );
  DFFPOSX1 arr_reg_42__7_ ( .D(n8151), .CLK(clk), .Q(arr[1393]) );
  DFFPOSX1 arr_reg_42__6_ ( .D(n8150), .CLK(clk), .Q(arr[1392]) );
  DFFPOSX1 arr_reg_42__5_ ( .D(n8149), .CLK(clk), .Q(arr[1391]) );
  DFFPOSX1 arr_reg_42__4_ ( .D(n8148), .CLK(clk), .Q(arr[1390]) );
  DFFPOSX1 arr_reg_42__3_ ( .D(n8147), .CLK(clk), .Q(arr[1389]) );
  DFFPOSX1 arr_reg_42__2_ ( .D(n8146), .CLK(clk), .Q(arr[1388]) );
  DFFPOSX1 arr_reg_42__1_ ( .D(n8145), .CLK(clk), .Q(arr[1387]) );
  DFFPOSX1 arr_reg_42__0_ ( .D(n8144), .CLK(clk), .Q(arr[1386]) );
  DFFPOSX1 arr_reg_41__32_ ( .D(n8143), .CLK(clk), .Q(arr[1385]) );
  DFFPOSX1 arr_reg_41__31_ ( .D(n8142), .CLK(clk), .Q(arr[1384]) );
  DFFPOSX1 arr_reg_41__30_ ( .D(n8141), .CLK(clk), .Q(arr[1383]) );
  DFFPOSX1 arr_reg_41__29_ ( .D(n8140), .CLK(clk), .Q(arr[1382]) );
  DFFPOSX1 arr_reg_41__28_ ( .D(n8139), .CLK(clk), .Q(arr[1381]) );
  DFFPOSX1 arr_reg_41__27_ ( .D(n8138), .CLK(clk), .Q(arr[1380]) );
  DFFPOSX1 arr_reg_41__26_ ( .D(n8137), .CLK(clk), .Q(arr[1379]) );
  DFFPOSX1 arr_reg_41__25_ ( .D(n8136), .CLK(clk), .Q(arr[1378]) );
  DFFPOSX1 arr_reg_41__24_ ( .D(n8135), .CLK(clk), .Q(arr[1377]) );
  DFFPOSX1 arr_reg_41__23_ ( .D(n8134), .CLK(clk), .Q(arr[1376]) );
  DFFPOSX1 arr_reg_41__22_ ( .D(n8133), .CLK(clk), .Q(arr[1375]) );
  DFFPOSX1 arr_reg_41__21_ ( .D(n8132), .CLK(clk), .Q(arr[1374]) );
  DFFPOSX1 arr_reg_41__20_ ( .D(n8131), .CLK(clk), .Q(arr[1373]) );
  DFFPOSX1 arr_reg_41__19_ ( .D(n8130), .CLK(clk), .Q(arr[1372]) );
  DFFPOSX1 arr_reg_41__18_ ( .D(n8129), .CLK(clk), .Q(arr[1371]) );
  DFFPOSX1 arr_reg_41__17_ ( .D(n8128), .CLK(clk), .Q(arr[1370]) );
  DFFPOSX1 arr_reg_41__16_ ( .D(n8127), .CLK(clk), .Q(arr[1369]) );
  DFFPOSX1 arr_reg_41__15_ ( .D(n8126), .CLK(clk), .Q(arr[1368]) );
  DFFPOSX1 arr_reg_41__14_ ( .D(n8125), .CLK(clk), .Q(arr[1367]) );
  DFFPOSX1 arr_reg_41__13_ ( .D(n8124), .CLK(clk), .Q(arr[1366]) );
  DFFPOSX1 arr_reg_41__12_ ( .D(n8123), .CLK(clk), .Q(arr[1365]) );
  DFFPOSX1 arr_reg_41__11_ ( .D(n8122), .CLK(clk), .Q(arr[1364]) );
  DFFPOSX1 arr_reg_41__10_ ( .D(n8121), .CLK(clk), .Q(arr[1363]) );
  DFFPOSX1 arr_reg_41__9_ ( .D(n8120), .CLK(clk), .Q(arr[1362]) );
  DFFPOSX1 arr_reg_41__8_ ( .D(n8119), .CLK(clk), .Q(arr[1361]) );
  DFFPOSX1 arr_reg_41__7_ ( .D(n8118), .CLK(clk), .Q(arr[1360]) );
  DFFPOSX1 arr_reg_41__6_ ( .D(n8117), .CLK(clk), .Q(arr[1359]) );
  DFFPOSX1 arr_reg_41__5_ ( .D(n8116), .CLK(clk), .Q(arr[1358]) );
  DFFPOSX1 arr_reg_41__4_ ( .D(n8115), .CLK(clk), .Q(arr[1357]) );
  DFFPOSX1 arr_reg_41__3_ ( .D(n8114), .CLK(clk), .Q(arr[1356]) );
  DFFPOSX1 arr_reg_41__2_ ( .D(n8113), .CLK(clk), .Q(arr[1355]) );
  DFFPOSX1 arr_reg_41__1_ ( .D(n8112), .CLK(clk), .Q(arr[1354]) );
  DFFPOSX1 arr_reg_41__0_ ( .D(n8111), .CLK(clk), .Q(arr[1353]) );
  DFFPOSX1 arr_reg_40__32_ ( .D(n8110), .CLK(clk), .Q(arr[1352]) );
  DFFPOSX1 arr_reg_40__31_ ( .D(n8109), .CLK(clk), .Q(arr[1351]) );
  DFFPOSX1 arr_reg_40__30_ ( .D(n8108), .CLK(clk), .Q(arr[1350]) );
  DFFPOSX1 arr_reg_40__29_ ( .D(n8107), .CLK(clk), .Q(arr[1349]) );
  DFFPOSX1 arr_reg_40__28_ ( .D(n8106), .CLK(clk), .Q(arr[1348]) );
  DFFPOSX1 arr_reg_40__27_ ( .D(n8105), .CLK(clk), .Q(arr[1347]) );
  DFFPOSX1 arr_reg_40__26_ ( .D(n8104), .CLK(clk), .Q(arr[1346]) );
  DFFPOSX1 arr_reg_40__25_ ( .D(n8103), .CLK(clk), .Q(arr[1345]) );
  DFFPOSX1 arr_reg_40__24_ ( .D(n8102), .CLK(clk), .Q(arr[1344]) );
  DFFPOSX1 arr_reg_40__23_ ( .D(n8101), .CLK(clk), .Q(arr[1343]) );
  DFFPOSX1 arr_reg_40__22_ ( .D(n8100), .CLK(clk), .Q(arr[1342]) );
  DFFPOSX1 arr_reg_40__21_ ( .D(n8099), .CLK(clk), .Q(arr[1341]) );
  DFFPOSX1 arr_reg_40__20_ ( .D(n8098), .CLK(clk), .Q(arr[1340]) );
  DFFPOSX1 arr_reg_40__19_ ( .D(n8097), .CLK(clk), .Q(arr[1339]) );
  DFFPOSX1 arr_reg_40__18_ ( .D(n8096), .CLK(clk), .Q(arr[1338]) );
  DFFPOSX1 arr_reg_40__17_ ( .D(n8095), .CLK(clk), .Q(arr[1337]) );
  DFFPOSX1 arr_reg_40__16_ ( .D(n8094), .CLK(clk), .Q(arr[1336]) );
  DFFPOSX1 arr_reg_40__15_ ( .D(n8093), .CLK(clk), .Q(arr[1335]) );
  DFFPOSX1 arr_reg_40__14_ ( .D(n8092), .CLK(clk), .Q(arr[1334]) );
  DFFPOSX1 arr_reg_40__13_ ( .D(n8091), .CLK(clk), .Q(arr[1333]) );
  DFFPOSX1 arr_reg_40__12_ ( .D(n8090), .CLK(clk), .Q(arr[1332]) );
  DFFPOSX1 arr_reg_40__11_ ( .D(n8089), .CLK(clk), .Q(arr[1331]) );
  DFFPOSX1 arr_reg_40__10_ ( .D(n8088), .CLK(clk), .Q(arr[1330]) );
  DFFPOSX1 arr_reg_40__9_ ( .D(n8087), .CLK(clk), .Q(arr[1329]) );
  DFFPOSX1 arr_reg_40__8_ ( .D(n8086), .CLK(clk), .Q(arr[1328]) );
  DFFPOSX1 arr_reg_40__7_ ( .D(n8085), .CLK(clk), .Q(arr[1327]) );
  DFFPOSX1 arr_reg_40__6_ ( .D(n8084), .CLK(clk), .Q(arr[1326]) );
  DFFPOSX1 arr_reg_40__5_ ( .D(n8083), .CLK(clk), .Q(arr[1325]) );
  DFFPOSX1 arr_reg_40__4_ ( .D(n8082), .CLK(clk), .Q(arr[1324]) );
  DFFPOSX1 arr_reg_40__3_ ( .D(n8081), .CLK(clk), .Q(arr[1323]) );
  DFFPOSX1 arr_reg_40__2_ ( .D(n8080), .CLK(clk), .Q(arr[1322]) );
  DFFPOSX1 arr_reg_40__1_ ( .D(n8079), .CLK(clk), .Q(arr[1321]) );
  DFFPOSX1 arr_reg_40__0_ ( .D(n8078), .CLK(clk), .Q(arr[1320]) );
  DFFPOSX1 arr_reg_39__32_ ( .D(n8077), .CLK(clk), .Q(arr[1319]) );
  DFFPOSX1 arr_reg_39__31_ ( .D(n8076), .CLK(clk), .Q(arr[1318]) );
  DFFPOSX1 arr_reg_39__30_ ( .D(n8075), .CLK(clk), .Q(arr[1317]) );
  DFFPOSX1 arr_reg_39__29_ ( .D(n8074), .CLK(clk), .Q(arr[1316]) );
  DFFPOSX1 arr_reg_39__28_ ( .D(n8073), .CLK(clk), .Q(arr[1315]) );
  DFFPOSX1 arr_reg_39__27_ ( .D(n8072), .CLK(clk), .Q(arr[1314]) );
  DFFPOSX1 arr_reg_39__26_ ( .D(n8071), .CLK(clk), .Q(arr[1313]) );
  DFFPOSX1 arr_reg_39__25_ ( .D(n8070), .CLK(clk), .Q(arr[1312]) );
  DFFPOSX1 arr_reg_39__24_ ( .D(n8069), .CLK(clk), .Q(arr[1311]) );
  DFFPOSX1 arr_reg_39__23_ ( .D(n8068), .CLK(clk), .Q(arr[1310]) );
  DFFPOSX1 arr_reg_39__22_ ( .D(n8067), .CLK(clk), .Q(arr[1309]) );
  DFFPOSX1 arr_reg_39__21_ ( .D(n8066), .CLK(clk), .Q(arr[1308]) );
  DFFPOSX1 arr_reg_39__20_ ( .D(n8065), .CLK(clk), .Q(arr[1307]) );
  DFFPOSX1 arr_reg_39__19_ ( .D(n8064), .CLK(clk), .Q(arr[1306]) );
  DFFPOSX1 arr_reg_39__18_ ( .D(n8063), .CLK(clk), .Q(arr[1305]) );
  DFFPOSX1 arr_reg_39__17_ ( .D(n8062), .CLK(clk), .Q(arr[1304]) );
  DFFPOSX1 arr_reg_39__16_ ( .D(n8061), .CLK(clk), .Q(arr[1303]) );
  DFFPOSX1 arr_reg_39__15_ ( .D(n8060), .CLK(clk), .Q(arr[1302]) );
  DFFPOSX1 arr_reg_39__14_ ( .D(n8059), .CLK(clk), .Q(arr[1301]) );
  DFFPOSX1 arr_reg_39__13_ ( .D(n8058), .CLK(clk), .Q(arr[1300]) );
  DFFPOSX1 arr_reg_39__12_ ( .D(n8057), .CLK(clk), .Q(arr[1299]) );
  DFFPOSX1 arr_reg_39__11_ ( .D(n8056), .CLK(clk), .Q(arr[1298]) );
  DFFPOSX1 arr_reg_39__10_ ( .D(n8055), .CLK(clk), .Q(arr[1297]) );
  DFFPOSX1 arr_reg_39__9_ ( .D(n8054), .CLK(clk), .Q(arr[1296]) );
  DFFPOSX1 arr_reg_39__8_ ( .D(n8053), .CLK(clk), .Q(arr[1295]) );
  DFFPOSX1 arr_reg_39__7_ ( .D(n8052), .CLK(clk), .Q(arr[1294]) );
  DFFPOSX1 arr_reg_39__6_ ( .D(n8051), .CLK(clk), .Q(arr[1293]) );
  DFFPOSX1 arr_reg_39__5_ ( .D(n8050), .CLK(clk), .Q(arr[1292]) );
  DFFPOSX1 arr_reg_39__4_ ( .D(n8049), .CLK(clk), .Q(arr[1291]) );
  DFFPOSX1 arr_reg_39__3_ ( .D(n8048), .CLK(clk), .Q(arr[1290]) );
  DFFPOSX1 arr_reg_39__2_ ( .D(n8047), .CLK(clk), .Q(arr[1289]) );
  DFFPOSX1 arr_reg_39__1_ ( .D(n8046), .CLK(clk), .Q(arr[1288]) );
  DFFPOSX1 arr_reg_39__0_ ( .D(n8045), .CLK(clk), .Q(arr[1287]) );
  DFFPOSX1 arr_reg_38__32_ ( .D(n8044), .CLK(clk), .Q(arr[1286]) );
  DFFPOSX1 arr_reg_38__31_ ( .D(n8043), .CLK(clk), .Q(arr[1285]) );
  DFFPOSX1 arr_reg_38__30_ ( .D(n8042), .CLK(clk), .Q(arr[1284]) );
  DFFPOSX1 arr_reg_38__29_ ( .D(n8041), .CLK(clk), .Q(arr[1283]) );
  DFFPOSX1 arr_reg_38__28_ ( .D(n8040), .CLK(clk), .Q(arr[1282]) );
  DFFPOSX1 arr_reg_38__27_ ( .D(n8039), .CLK(clk), .Q(arr[1281]) );
  DFFPOSX1 arr_reg_38__26_ ( .D(n8038), .CLK(clk), .Q(arr[1280]) );
  DFFPOSX1 arr_reg_38__25_ ( .D(n8037), .CLK(clk), .Q(arr[1279]) );
  DFFPOSX1 arr_reg_38__24_ ( .D(n8036), .CLK(clk), .Q(arr[1278]) );
  DFFPOSX1 arr_reg_38__23_ ( .D(n8035), .CLK(clk), .Q(arr[1277]) );
  DFFPOSX1 arr_reg_38__22_ ( .D(n8034), .CLK(clk), .Q(arr[1276]) );
  DFFPOSX1 arr_reg_38__21_ ( .D(n8033), .CLK(clk), .Q(arr[1275]) );
  DFFPOSX1 arr_reg_38__20_ ( .D(n8032), .CLK(clk), .Q(arr[1274]) );
  DFFPOSX1 arr_reg_38__19_ ( .D(n8031), .CLK(clk), .Q(arr[1273]) );
  DFFPOSX1 arr_reg_38__18_ ( .D(n8030), .CLK(clk), .Q(arr[1272]) );
  DFFPOSX1 arr_reg_38__17_ ( .D(n8029), .CLK(clk), .Q(arr[1271]) );
  DFFPOSX1 arr_reg_38__16_ ( .D(n8028), .CLK(clk), .Q(arr[1270]) );
  DFFPOSX1 arr_reg_38__15_ ( .D(n8027), .CLK(clk), .Q(arr[1269]) );
  DFFPOSX1 arr_reg_38__14_ ( .D(n8026), .CLK(clk), .Q(arr[1268]) );
  DFFPOSX1 arr_reg_38__13_ ( .D(n8025), .CLK(clk), .Q(arr[1267]) );
  DFFPOSX1 arr_reg_38__12_ ( .D(n8024), .CLK(clk), .Q(arr[1266]) );
  DFFPOSX1 arr_reg_38__11_ ( .D(n8023), .CLK(clk), .Q(arr[1265]) );
  DFFPOSX1 arr_reg_38__10_ ( .D(n8022), .CLK(clk), .Q(arr[1264]) );
  DFFPOSX1 arr_reg_38__9_ ( .D(n8021), .CLK(clk), .Q(arr[1263]) );
  DFFPOSX1 arr_reg_38__8_ ( .D(n8020), .CLK(clk), .Q(arr[1262]) );
  DFFPOSX1 arr_reg_38__7_ ( .D(n8019), .CLK(clk), .Q(arr[1261]) );
  DFFPOSX1 arr_reg_38__6_ ( .D(n8018), .CLK(clk), .Q(arr[1260]) );
  DFFPOSX1 arr_reg_38__5_ ( .D(n8017), .CLK(clk), .Q(arr[1259]) );
  DFFPOSX1 arr_reg_38__4_ ( .D(n8016), .CLK(clk), .Q(arr[1258]) );
  DFFPOSX1 arr_reg_38__3_ ( .D(n8015), .CLK(clk), .Q(arr[1257]) );
  DFFPOSX1 arr_reg_38__2_ ( .D(n8014), .CLK(clk), .Q(arr[1256]) );
  DFFPOSX1 arr_reg_38__1_ ( .D(n8013), .CLK(clk), .Q(arr[1255]) );
  DFFPOSX1 arr_reg_38__0_ ( .D(n8012), .CLK(clk), .Q(arr[1254]) );
  DFFPOSX1 arr_reg_37__32_ ( .D(n8011), .CLK(clk), .Q(arr[1253]) );
  DFFPOSX1 arr_reg_37__31_ ( .D(n8010), .CLK(clk), .Q(arr[1252]) );
  DFFPOSX1 arr_reg_37__30_ ( .D(n8009), .CLK(clk), .Q(arr[1251]) );
  DFFPOSX1 arr_reg_37__29_ ( .D(n8008), .CLK(clk), .Q(arr[1250]) );
  DFFPOSX1 arr_reg_37__28_ ( .D(n8007), .CLK(clk), .Q(arr[1249]) );
  DFFPOSX1 arr_reg_37__27_ ( .D(n8006), .CLK(clk), .Q(arr[1248]) );
  DFFPOSX1 arr_reg_37__26_ ( .D(n8005), .CLK(clk), .Q(arr[1247]) );
  DFFPOSX1 arr_reg_37__25_ ( .D(n8004), .CLK(clk), .Q(arr[1246]) );
  DFFPOSX1 arr_reg_37__24_ ( .D(n8003), .CLK(clk), .Q(arr[1245]) );
  DFFPOSX1 arr_reg_37__23_ ( .D(n8002), .CLK(clk), .Q(arr[1244]) );
  DFFPOSX1 arr_reg_37__22_ ( .D(n8001), .CLK(clk), .Q(arr[1243]) );
  DFFPOSX1 arr_reg_37__21_ ( .D(n8000), .CLK(clk), .Q(arr[1242]) );
  DFFPOSX1 arr_reg_37__20_ ( .D(n7999), .CLK(clk), .Q(arr[1241]) );
  DFFPOSX1 arr_reg_37__19_ ( .D(n7998), .CLK(clk), .Q(arr[1240]) );
  DFFPOSX1 arr_reg_37__18_ ( .D(n7997), .CLK(clk), .Q(arr[1239]) );
  DFFPOSX1 arr_reg_37__17_ ( .D(n7996), .CLK(clk), .Q(arr[1238]) );
  DFFPOSX1 arr_reg_37__16_ ( .D(n7995), .CLK(clk), .Q(arr[1237]) );
  DFFPOSX1 arr_reg_37__15_ ( .D(n7994), .CLK(clk), .Q(arr[1236]) );
  DFFPOSX1 arr_reg_37__14_ ( .D(n7993), .CLK(clk), .Q(arr[1235]) );
  DFFPOSX1 arr_reg_37__13_ ( .D(n7992), .CLK(clk), .Q(arr[1234]) );
  DFFPOSX1 arr_reg_37__12_ ( .D(n7991), .CLK(clk), .Q(arr[1233]) );
  DFFPOSX1 arr_reg_37__11_ ( .D(n7990), .CLK(clk), .Q(arr[1232]) );
  DFFPOSX1 arr_reg_37__10_ ( .D(n7989), .CLK(clk), .Q(arr[1231]) );
  DFFPOSX1 arr_reg_37__9_ ( .D(n7988), .CLK(clk), .Q(arr[1230]) );
  DFFPOSX1 arr_reg_37__8_ ( .D(n7987), .CLK(clk), .Q(arr[1229]) );
  DFFPOSX1 arr_reg_37__7_ ( .D(n7986), .CLK(clk), .Q(arr[1228]) );
  DFFPOSX1 arr_reg_37__6_ ( .D(n7985), .CLK(clk), .Q(arr[1227]) );
  DFFPOSX1 arr_reg_37__5_ ( .D(n7984), .CLK(clk), .Q(arr[1226]) );
  DFFPOSX1 arr_reg_37__4_ ( .D(n7983), .CLK(clk), .Q(arr[1225]) );
  DFFPOSX1 arr_reg_37__3_ ( .D(n7982), .CLK(clk), .Q(arr[1224]) );
  DFFPOSX1 arr_reg_37__2_ ( .D(n7981), .CLK(clk), .Q(arr[1223]) );
  DFFPOSX1 arr_reg_37__1_ ( .D(n7980), .CLK(clk), .Q(arr[1222]) );
  DFFPOSX1 arr_reg_37__0_ ( .D(n7979), .CLK(clk), .Q(arr[1221]) );
  DFFPOSX1 arr_reg_36__32_ ( .D(n7978), .CLK(clk), .Q(arr[1220]) );
  DFFPOSX1 arr_reg_36__31_ ( .D(n7977), .CLK(clk), .Q(arr[1219]) );
  DFFPOSX1 arr_reg_36__30_ ( .D(n7976), .CLK(clk), .Q(arr[1218]) );
  DFFPOSX1 arr_reg_36__29_ ( .D(n7975), .CLK(clk), .Q(arr[1217]) );
  DFFPOSX1 arr_reg_36__28_ ( .D(n7974), .CLK(clk), .Q(arr[1216]) );
  DFFPOSX1 arr_reg_36__27_ ( .D(n7973), .CLK(clk), .Q(arr[1215]) );
  DFFPOSX1 arr_reg_36__26_ ( .D(n7972), .CLK(clk), .Q(arr[1214]) );
  DFFPOSX1 arr_reg_36__25_ ( .D(n7971), .CLK(clk), .Q(arr[1213]) );
  DFFPOSX1 arr_reg_36__24_ ( .D(n7970), .CLK(clk), .Q(arr[1212]) );
  DFFPOSX1 arr_reg_36__23_ ( .D(n7969), .CLK(clk), .Q(arr[1211]) );
  DFFPOSX1 arr_reg_36__22_ ( .D(n7968), .CLK(clk), .Q(arr[1210]) );
  DFFPOSX1 arr_reg_36__21_ ( .D(n7967), .CLK(clk), .Q(arr[1209]) );
  DFFPOSX1 arr_reg_36__20_ ( .D(n7966), .CLK(clk), .Q(arr[1208]) );
  DFFPOSX1 arr_reg_36__19_ ( .D(n7965), .CLK(clk), .Q(arr[1207]) );
  DFFPOSX1 arr_reg_36__18_ ( .D(n7964), .CLK(clk), .Q(arr[1206]) );
  DFFPOSX1 arr_reg_36__17_ ( .D(n7963), .CLK(clk), .Q(arr[1205]) );
  DFFPOSX1 arr_reg_36__16_ ( .D(n7962), .CLK(clk), .Q(arr[1204]) );
  DFFPOSX1 arr_reg_36__15_ ( .D(n7961), .CLK(clk), .Q(arr[1203]) );
  DFFPOSX1 arr_reg_36__14_ ( .D(n7960), .CLK(clk), .Q(arr[1202]) );
  DFFPOSX1 arr_reg_36__13_ ( .D(n7959), .CLK(clk), .Q(arr[1201]) );
  DFFPOSX1 arr_reg_36__12_ ( .D(n7958), .CLK(clk), .Q(arr[1200]) );
  DFFPOSX1 arr_reg_36__11_ ( .D(n7957), .CLK(clk), .Q(arr[1199]) );
  DFFPOSX1 arr_reg_36__10_ ( .D(n7956), .CLK(clk), .Q(arr[1198]) );
  DFFPOSX1 arr_reg_36__9_ ( .D(n7955), .CLK(clk), .Q(arr[1197]) );
  DFFPOSX1 arr_reg_36__8_ ( .D(n7954), .CLK(clk), .Q(arr[1196]) );
  DFFPOSX1 arr_reg_36__7_ ( .D(n7953), .CLK(clk), .Q(arr[1195]) );
  DFFPOSX1 arr_reg_36__6_ ( .D(n7952), .CLK(clk), .Q(arr[1194]) );
  DFFPOSX1 arr_reg_36__5_ ( .D(n7951), .CLK(clk), .Q(arr[1193]) );
  DFFPOSX1 arr_reg_36__4_ ( .D(n7950), .CLK(clk), .Q(arr[1192]) );
  DFFPOSX1 arr_reg_36__3_ ( .D(n7949), .CLK(clk), .Q(arr[1191]) );
  DFFPOSX1 arr_reg_36__2_ ( .D(n7948), .CLK(clk), .Q(arr[1190]) );
  DFFPOSX1 arr_reg_36__1_ ( .D(n7947), .CLK(clk), .Q(arr[1189]) );
  DFFPOSX1 arr_reg_36__0_ ( .D(n7946), .CLK(clk), .Q(arr[1188]) );
  DFFPOSX1 arr_reg_35__32_ ( .D(n7945), .CLK(clk), .Q(arr[1187]) );
  DFFPOSX1 arr_reg_35__31_ ( .D(n7944), .CLK(clk), .Q(arr[1186]) );
  DFFPOSX1 arr_reg_35__30_ ( .D(n7943), .CLK(clk), .Q(arr[1185]) );
  DFFPOSX1 arr_reg_35__29_ ( .D(n7942), .CLK(clk), .Q(arr[1184]) );
  DFFPOSX1 arr_reg_35__28_ ( .D(n7941), .CLK(clk), .Q(arr[1183]) );
  DFFPOSX1 arr_reg_35__27_ ( .D(n7940), .CLK(clk), .Q(arr[1182]) );
  DFFPOSX1 arr_reg_35__26_ ( .D(n7939), .CLK(clk), .Q(arr[1181]) );
  DFFPOSX1 arr_reg_35__25_ ( .D(n7938), .CLK(clk), .Q(arr[1180]) );
  DFFPOSX1 arr_reg_35__24_ ( .D(n7937), .CLK(clk), .Q(arr[1179]) );
  DFFPOSX1 arr_reg_35__23_ ( .D(n7936), .CLK(clk), .Q(arr[1178]) );
  DFFPOSX1 arr_reg_35__22_ ( .D(n7935), .CLK(clk), .Q(arr[1177]) );
  DFFPOSX1 arr_reg_35__21_ ( .D(n7934), .CLK(clk), .Q(arr[1176]) );
  DFFPOSX1 arr_reg_35__20_ ( .D(n7933), .CLK(clk), .Q(arr[1175]) );
  DFFPOSX1 arr_reg_35__19_ ( .D(n7932), .CLK(clk), .Q(arr[1174]) );
  DFFPOSX1 arr_reg_35__18_ ( .D(n7931), .CLK(clk), .Q(arr[1173]) );
  DFFPOSX1 arr_reg_35__17_ ( .D(n7930), .CLK(clk), .Q(arr[1172]) );
  DFFPOSX1 arr_reg_35__16_ ( .D(n7929), .CLK(clk), .Q(arr[1171]) );
  DFFPOSX1 arr_reg_35__15_ ( .D(n7928), .CLK(clk), .Q(arr[1170]) );
  DFFPOSX1 arr_reg_35__14_ ( .D(n7927), .CLK(clk), .Q(arr[1169]) );
  DFFPOSX1 arr_reg_35__13_ ( .D(n7926), .CLK(clk), .Q(arr[1168]) );
  DFFPOSX1 arr_reg_35__12_ ( .D(n7925), .CLK(clk), .Q(arr[1167]) );
  DFFPOSX1 arr_reg_35__11_ ( .D(n7924), .CLK(clk), .Q(arr[1166]) );
  DFFPOSX1 arr_reg_35__10_ ( .D(n7923), .CLK(clk), .Q(arr[1165]) );
  DFFPOSX1 arr_reg_35__9_ ( .D(n7922), .CLK(clk), .Q(arr[1164]) );
  DFFPOSX1 arr_reg_35__8_ ( .D(n7921), .CLK(clk), .Q(arr[1163]) );
  DFFPOSX1 arr_reg_35__7_ ( .D(n7920), .CLK(clk), .Q(arr[1162]) );
  DFFPOSX1 arr_reg_35__6_ ( .D(n7919), .CLK(clk), .Q(arr[1161]) );
  DFFPOSX1 arr_reg_35__5_ ( .D(n7918), .CLK(clk), .Q(arr[1160]) );
  DFFPOSX1 arr_reg_35__4_ ( .D(n7917), .CLK(clk), .Q(arr[1159]) );
  DFFPOSX1 arr_reg_35__3_ ( .D(n7916), .CLK(clk), .Q(arr[1158]) );
  DFFPOSX1 arr_reg_35__2_ ( .D(n7915), .CLK(clk), .Q(arr[1157]) );
  DFFPOSX1 arr_reg_35__1_ ( .D(n7914), .CLK(clk), .Q(arr[1156]) );
  DFFPOSX1 arr_reg_35__0_ ( .D(n7913), .CLK(clk), .Q(arr[1155]) );
  DFFPOSX1 arr_reg_34__32_ ( .D(n7912), .CLK(clk), .Q(arr[1154]) );
  DFFPOSX1 arr_reg_34__31_ ( .D(n7911), .CLK(clk), .Q(arr[1153]) );
  DFFPOSX1 arr_reg_34__30_ ( .D(n7910), .CLK(clk), .Q(arr[1152]) );
  DFFPOSX1 arr_reg_34__29_ ( .D(n7909), .CLK(clk), .Q(arr[1151]) );
  DFFPOSX1 arr_reg_34__28_ ( .D(n7908), .CLK(clk), .Q(arr[1150]) );
  DFFPOSX1 arr_reg_34__27_ ( .D(n7907), .CLK(clk), .Q(arr[1149]) );
  DFFPOSX1 arr_reg_34__26_ ( .D(n7906), .CLK(clk), .Q(arr[1148]) );
  DFFPOSX1 arr_reg_34__25_ ( .D(n7905), .CLK(clk), .Q(arr[1147]) );
  DFFPOSX1 arr_reg_34__24_ ( .D(n7904), .CLK(clk), .Q(arr[1146]) );
  DFFPOSX1 arr_reg_34__23_ ( .D(n7903), .CLK(clk), .Q(arr[1145]) );
  DFFPOSX1 arr_reg_34__22_ ( .D(n7902), .CLK(clk), .Q(arr[1144]) );
  DFFPOSX1 arr_reg_34__21_ ( .D(n7901), .CLK(clk), .Q(arr[1143]) );
  DFFPOSX1 arr_reg_34__20_ ( .D(n7900), .CLK(clk), .Q(arr[1142]) );
  DFFPOSX1 arr_reg_34__19_ ( .D(n7899), .CLK(clk), .Q(arr[1141]) );
  DFFPOSX1 arr_reg_34__18_ ( .D(n7898), .CLK(clk), .Q(arr[1140]) );
  DFFPOSX1 arr_reg_34__17_ ( .D(n7897), .CLK(clk), .Q(arr[1139]) );
  DFFPOSX1 arr_reg_34__16_ ( .D(n7896), .CLK(clk), .Q(arr[1138]) );
  DFFPOSX1 arr_reg_34__15_ ( .D(n7895), .CLK(clk), .Q(arr[1137]) );
  DFFPOSX1 arr_reg_34__14_ ( .D(n7894), .CLK(clk), .Q(arr[1136]) );
  DFFPOSX1 arr_reg_34__13_ ( .D(n7893), .CLK(clk), .Q(arr[1135]) );
  DFFPOSX1 arr_reg_34__12_ ( .D(n7892), .CLK(clk), .Q(arr[1134]) );
  DFFPOSX1 arr_reg_34__11_ ( .D(n7891), .CLK(clk), .Q(arr[1133]) );
  DFFPOSX1 arr_reg_34__10_ ( .D(n7890), .CLK(clk), .Q(arr[1132]) );
  DFFPOSX1 arr_reg_34__9_ ( .D(n7889), .CLK(clk), .Q(arr[1131]) );
  DFFPOSX1 arr_reg_34__8_ ( .D(n7888), .CLK(clk), .Q(arr[1130]) );
  DFFPOSX1 arr_reg_34__7_ ( .D(n7887), .CLK(clk), .Q(arr[1129]) );
  DFFPOSX1 arr_reg_34__6_ ( .D(n7886), .CLK(clk), .Q(arr[1128]) );
  DFFPOSX1 arr_reg_34__5_ ( .D(n7885), .CLK(clk), .Q(arr[1127]) );
  DFFPOSX1 arr_reg_34__4_ ( .D(n7884), .CLK(clk), .Q(arr[1126]) );
  DFFPOSX1 arr_reg_34__3_ ( .D(n7883), .CLK(clk), .Q(arr[1125]) );
  DFFPOSX1 arr_reg_34__2_ ( .D(n7882), .CLK(clk), .Q(arr[1124]) );
  DFFPOSX1 arr_reg_34__1_ ( .D(n7881), .CLK(clk), .Q(arr[1123]) );
  DFFPOSX1 arr_reg_34__0_ ( .D(n7880), .CLK(clk), .Q(arr[1122]) );
  DFFPOSX1 arr_reg_33__32_ ( .D(n7879), .CLK(clk), .Q(arr[1121]) );
  DFFPOSX1 arr_reg_33__31_ ( .D(n7878), .CLK(clk), .Q(arr[1120]) );
  DFFPOSX1 arr_reg_33__30_ ( .D(n7877), .CLK(clk), .Q(arr[1119]) );
  DFFPOSX1 arr_reg_33__29_ ( .D(n7876), .CLK(clk), .Q(arr[1118]) );
  DFFPOSX1 arr_reg_33__28_ ( .D(n7875), .CLK(clk), .Q(arr[1117]) );
  DFFPOSX1 arr_reg_33__27_ ( .D(n7874), .CLK(clk), .Q(arr[1116]) );
  DFFPOSX1 arr_reg_33__26_ ( .D(n7873), .CLK(clk), .Q(arr[1115]) );
  DFFPOSX1 arr_reg_33__25_ ( .D(n7872), .CLK(clk), .Q(arr[1114]) );
  DFFPOSX1 arr_reg_33__24_ ( .D(n7871), .CLK(clk), .Q(arr[1113]) );
  DFFPOSX1 arr_reg_33__23_ ( .D(n7870), .CLK(clk), .Q(arr[1112]) );
  DFFPOSX1 arr_reg_33__22_ ( .D(n7869), .CLK(clk), .Q(arr[1111]) );
  DFFPOSX1 arr_reg_33__21_ ( .D(n7868), .CLK(clk), .Q(arr[1110]) );
  DFFPOSX1 arr_reg_33__20_ ( .D(n7867), .CLK(clk), .Q(arr[1109]) );
  DFFPOSX1 arr_reg_33__19_ ( .D(n7866), .CLK(clk), .Q(arr[1108]) );
  DFFPOSX1 arr_reg_33__18_ ( .D(n7865), .CLK(clk), .Q(arr[1107]) );
  DFFPOSX1 arr_reg_33__17_ ( .D(n7864), .CLK(clk), .Q(arr[1106]) );
  DFFPOSX1 arr_reg_33__16_ ( .D(n7863), .CLK(clk), .Q(arr[1105]) );
  DFFPOSX1 arr_reg_33__15_ ( .D(n7862), .CLK(clk), .Q(arr[1104]) );
  DFFPOSX1 arr_reg_33__14_ ( .D(n7861), .CLK(clk), .Q(arr[1103]) );
  DFFPOSX1 arr_reg_33__13_ ( .D(n7860), .CLK(clk), .Q(arr[1102]) );
  DFFPOSX1 arr_reg_33__12_ ( .D(n7859), .CLK(clk), .Q(arr[1101]) );
  DFFPOSX1 arr_reg_33__11_ ( .D(n7858), .CLK(clk), .Q(arr[1100]) );
  DFFPOSX1 arr_reg_33__10_ ( .D(n7857), .CLK(clk), .Q(arr[1099]) );
  DFFPOSX1 arr_reg_33__9_ ( .D(n7856), .CLK(clk), .Q(arr[1098]) );
  DFFPOSX1 arr_reg_33__8_ ( .D(n7855), .CLK(clk), .Q(arr[1097]) );
  DFFPOSX1 arr_reg_33__7_ ( .D(n7854), .CLK(clk), .Q(arr[1096]) );
  DFFPOSX1 arr_reg_33__6_ ( .D(n7853), .CLK(clk), .Q(arr[1095]) );
  DFFPOSX1 arr_reg_33__5_ ( .D(n7852), .CLK(clk), .Q(arr[1094]) );
  DFFPOSX1 arr_reg_33__4_ ( .D(n7851), .CLK(clk), .Q(arr[1093]) );
  DFFPOSX1 arr_reg_33__3_ ( .D(n7850), .CLK(clk), .Q(arr[1092]) );
  DFFPOSX1 arr_reg_33__2_ ( .D(n7849), .CLK(clk), .Q(arr[1091]) );
  DFFPOSX1 arr_reg_33__1_ ( .D(n7848), .CLK(clk), .Q(arr[1090]) );
  DFFPOSX1 arr_reg_33__0_ ( .D(n7847), .CLK(clk), .Q(arr[1089]) );
  DFFPOSX1 arr_reg_32__32_ ( .D(n7846), .CLK(clk), .Q(arr[1088]) );
  DFFPOSX1 arr_reg_32__31_ ( .D(n7845), .CLK(clk), .Q(arr[1087]) );
  DFFPOSX1 arr_reg_32__30_ ( .D(n7844), .CLK(clk), .Q(arr[1086]) );
  DFFPOSX1 arr_reg_32__29_ ( .D(n7843), .CLK(clk), .Q(arr[1085]) );
  DFFPOSX1 arr_reg_32__28_ ( .D(n7842), .CLK(clk), .Q(arr[1084]) );
  DFFPOSX1 arr_reg_32__27_ ( .D(n7841), .CLK(clk), .Q(arr[1083]) );
  DFFPOSX1 arr_reg_32__26_ ( .D(n7840), .CLK(clk), .Q(arr[1082]) );
  DFFPOSX1 arr_reg_32__25_ ( .D(n7839), .CLK(clk), .Q(arr[1081]) );
  DFFPOSX1 arr_reg_32__24_ ( .D(n7838), .CLK(clk), .Q(arr[1080]) );
  DFFPOSX1 arr_reg_32__23_ ( .D(n7837), .CLK(clk), .Q(arr[1079]) );
  DFFPOSX1 arr_reg_32__22_ ( .D(n7836), .CLK(clk), .Q(arr[1078]) );
  DFFPOSX1 arr_reg_32__21_ ( .D(n7835), .CLK(clk), .Q(arr[1077]) );
  DFFPOSX1 arr_reg_32__20_ ( .D(n7834), .CLK(clk), .Q(arr[1076]) );
  DFFPOSX1 arr_reg_32__19_ ( .D(n7833), .CLK(clk), .Q(arr[1075]) );
  DFFPOSX1 arr_reg_32__18_ ( .D(n7832), .CLK(clk), .Q(arr[1074]) );
  DFFPOSX1 arr_reg_32__17_ ( .D(n7831), .CLK(clk), .Q(arr[1073]) );
  DFFPOSX1 arr_reg_32__16_ ( .D(n7830), .CLK(clk), .Q(arr[1072]) );
  DFFPOSX1 arr_reg_32__15_ ( .D(n7829), .CLK(clk), .Q(arr[1071]) );
  DFFPOSX1 arr_reg_32__14_ ( .D(n7828), .CLK(clk), .Q(arr[1070]) );
  DFFPOSX1 arr_reg_32__13_ ( .D(n7827), .CLK(clk), .Q(arr[1069]) );
  DFFPOSX1 arr_reg_32__12_ ( .D(n7826), .CLK(clk), .Q(arr[1068]) );
  DFFPOSX1 arr_reg_32__11_ ( .D(n7825), .CLK(clk), .Q(arr[1067]) );
  DFFPOSX1 arr_reg_32__10_ ( .D(n7824), .CLK(clk), .Q(arr[1066]) );
  DFFPOSX1 arr_reg_32__9_ ( .D(n7823), .CLK(clk), .Q(arr[1065]) );
  DFFPOSX1 arr_reg_32__8_ ( .D(n7822), .CLK(clk), .Q(arr[1064]) );
  DFFPOSX1 arr_reg_32__7_ ( .D(n7821), .CLK(clk), .Q(arr[1063]) );
  DFFPOSX1 arr_reg_32__6_ ( .D(n7820), .CLK(clk), .Q(arr[1062]) );
  DFFPOSX1 arr_reg_32__5_ ( .D(n7819), .CLK(clk), .Q(arr[1061]) );
  DFFPOSX1 arr_reg_32__4_ ( .D(n7818), .CLK(clk), .Q(arr[1060]) );
  DFFPOSX1 arr_reg_32__3_ ( .D(n7817), .CLK(clk), .Q(arr[1059]) );
  DFFPOSX1 arr_reg_32__2_ ( .D(n7816), .CLK(clk), .Q(arr[1058]) );
  DFFPOSX1 arr_reg_32__1_ ( .D(n7815), .CLK(clk), .Q(arr[1057]) );
  DFFPOSX1 arr_reg_32__0_ ( .D(n7814), .CLK(clk), .Q(arr[1056]) );
  DFFPOSX1 arr_reg_31__32_ ( .D(n7813), .CLK(clk), .Q(arr[1055]) );
  DFFPOSX1 arr_reg_31__31_ ( .D(n7812), .CLK(clk), .Q(arr[1054]) );
  DFFPOSX1 arr_reg_31__30_ ( .D(n7811), .CLK(clk), .Q(arr[1053]) );
  DFFPOSX1 arr_reg_31__29_ ( .D(n7810), .CLK(clk), .Q(arr[1052]) );
  DFFPOSX1 arr_reg_31__28_ ( .D(n7809), .CLK(clk), .Q(arr[1051]) );
  DFFPOSX1 arr_reg_31__27_ ( .D(n7808), .CLK(clk), .Q(arr[1050]) );
  DFFPOSX1 arr_reg_31__26_ ( .D(n7807), .CLK(clk), .Q(arr[1049]) );
  DFFPOSX1 arr_reg_31__25_ ( .D(n7806), .CLK(clk), .Q(arr[1048]) );
  DFFPOSX1 arr_reg_31__24_ ( .D(n7805), .CLK(clk), .Q(arr[1047]) );
  DFFPOSX1 arr_reg_31__23_ ( .D(n7804), .CLK(clk), .Q(arr[1046]) );
  DFFPOSX1 arr_reg_31__22_ ( .D(n7803), .CLK(clk), .Q(arr[1045]) );
  DFFPOSX1 arr_reg_31__21_ ( .D(n7802), .CLK(clk), .Q(arr[1044]) );
  DFFPOSX1 arr_reg_31__20_ ( .D(n7801), .CLK(clk), .Q(arr[1043]) );
  DFFPOSX1 arr_reg_31__19_ ( .D(n7800), .CLK(clk), .Q(arr[1042]) );
  DFFPOSX1 arr_reg_31__18_ ( .D(n7799), .CLK(clk), .Q(arr[1041]) );
  DFFPOSX1 arr_reg_31__17_ ( .D(n7798), .CLK(clk), .Q(arr[1040]) );
  DFFPOSX1 arr_reg_31__16_ ( .D(n7797), .CLK(clk), .Q(arr[1039]) );
  DFFPOSX1 arr_reg_31__15_ ( .D(n7796), .CLK(clk), .Q(arr[1038]) );
  DFFPOSX1 arr_reg_31__14_ ( .D(n7795), .CLK(clk), .Q(arr[1037]) );
  DFFPOSX1 arr_reg_31__13_ ( .D(n7794), .CLK(clk), .Q(arr[1036]) );
  DFFPOSX1 arr_reg_31__12_ ( .D(n7793), .CLK(clk), .Q(arr[1035]) );
  DFFPOSX1 arr_reg_31__11_ ( .D(n7792), .CLK(clk), .Q(arr[1034]) );
  DFFPOSX1 arr_reg_31__10_ ( .D(n7791), .CLK(clk), .Q(arr[1033]) );
  DFFPOSX1 arr_reg_31__9_ ( .D(n7790), .CLK(clk), .Q(arr[1032]) );
  DFFPOSX1 arr_reg_31__8_ ( .D(n7789), .CLK(clk), .Q(arr[1031]) );
  DFFPOSX1 arr_reg_31__7_ ( .D(n7788), .CLK(clk), .Q(arr[1030]) );
  DFFPOSX1 arr_reg_31__6_ ( .D(n7787), .CLK(clk), .Q(arr[1029]) );
  DFFPOSX1 arr_reg_31__5_ ( .D(n7786), .CLK(clk), .Q(arr[1028]) );
  DFFPOSX1 arr_reg_31__4_ ( .D(n7785), .CLK(clk), .Q(arr[1027]) );
  DFFPOSX1 arr_reg_31__3_ ( .D(n7784), .CLK(clk), .Q(arr[1026]) );
  DFFPOSX1 arr_reg_31__2_ ( .D(n7783), .CLK(clk), .Q(arr[1025]) );
  DFFPOSX1 arr_reg_31__1_ ( .D(n7782), .CLK(clk), .Q(arr[1024]) );
  DFFPOSX1 arr_reg_31__0_ ( .D(n7781), .CLK(clk), .Q(arr[1023]) );
  DFFPOSX1 arr_reg_30__32_ ( .D(n7780), .CLK(clk), .Q(arr[1022]) );
  DFFPOSX1 arr_reg_30__31_ ( .D(n7779), .CLK(clk), .Q(arr[1021]) );
  DFFPOSX1 arr_reg_30__30_ ( .D(n7778), .CLK(clk), .Q(arr[1020]) );
  DFFPOSX1 arr_reg_30__29_ ( .D(n7777), .CLK(clk), .Q(arr[1019]) );
  DFFPOSX1 arr_reg_30__28_ ( .D(n7776), .CLK(clk), .Q(arr[1018]) );
  DFFPOSX1 arr_reg_30__27_ ( .D(n7775), .CLK(clk), .Q(arr[1017]) );
  DFFPOSX1 arr_reg_30__26_ ( .D(n7774), .CLK(clk), .Q(arr[1016]) );
  DFFPOSX1 arr_reg_30__25_ ( .D(n7773), .CLK(clk), .Q(arr[1015]) );
  DFFPOSX1 arr_reg_30__24_ ( .D(n7772), .CLK(clk), .Q(arr[1014]) );
  DFFPOSX1 arr_reg_30__23_ ( .D(n7771), .CLK(clk), .Q(arr[1013]) );
  DFFPOSX1 arr_reg_30__22_ ( .D(n7770), .CLK(clk), .Q(arr[1012]) );
  DFFPOSX1 arr_reg_30__21_ ( .D(n7769), .CLK(clk), .Q(arr[1011]) );
  DFFPOSX1 arr_reg_30__20_ ( .D(n7768), .CLK(clk), .Q(arr[1010]) );
  DFFPOSX1 arr_reg_30__19_ ( .D(n7767), .CLK(clk), .Q(arr[1009]) );
  DFFPOSX1 arr_reg_30__18_ ( .D(n7766), .CLK(clk), .Q(arr[1008]) );
  DFFPOSX1 arr_reg_30__17_ ( .D(n7765), .CLK(clk), .Q(arr[1007]) );
  DFFPOSX1 arr_reg_30__16_ ( .D(n7764), .CLK(clk), .Q(arr[1006]) );
  DFFPOSX1 arr_reg_30__15_ ( .D(n7763), .CLK(clk), .Q(arr[1005]) );
  DFFPOSX1 arr_reg_30__14_ ( .D(n7762), .CLK(clk), .Q(arr[1004]) );
  DFFPOSX1 arr_reg_30__13_ ( .D(n7761), .CLK(clk), .Q(arr[1003]) );
  DFFPOSX1 arr_reg_30__12_ ( .D(n7760), .CLK(clk), .Q(arr[1002]) );
  DFFPOSX1 arr_reg_30__11_ ( .D(n7759), .CLK(clk), .Q(arr[1001]) );
  DFFPOSX1 arr_reg_30__10_ ( .D(n7758), .CLK(clk), .Q(arr[1000]) );
  DFFPOSX1 arr_reg_30__9_ ( .D(n7757), .CLK(clk), .Q(arr[999]) );
  DFFPOSX1 arr_reg_30__8_ ( .D(n7756), .CLK(clk), .Q(arr[998]) );
  DFFPOSX1 arr_reg_30__7_ ( .D(n7755), .CLK(clk), .Q(arr[997]) );
  DFFPOSX1 arr_reg_30__6_ ( .D(n7754), .CLK(clk), .Q(arr[996]) );
  DFFPOSX1 arr_reg_30__5_ ( .D(n7753), .CLK(clk), .Q(arr[995]) );
  DFFPOSX1 arr_reg_30__4_ ( .D(n7752), .CLK(clk), .Q(arr[994]) );
  DFFPOSX1 arr_reg_30__3_ ( .D(n7751), .CLK(clk), .Q(arr[993]) );
  DFFPOSX1 arr_reg_30__2_ ( .D(n7750), .CLK(clk), .Q(arr[992]) );
  DFFPOSX1 arr_reg_30__1_ ( .D(n7749), .CLK(clk), .Q(arr[991]) );
  DFFPOSX1 arr_reg_30__0_ ( .D(n7748), .CLK(clk), .Q(arr[990]) );
  DFFPOSX1 arr_reg_29__32_ ( .D(n7747), .CLK(clk), .Q(arr[989]) );
  DFFPOSX1 arr_reg_29__31_ ( .D(n7746), .CLK(clk), .Q(arr[988]) );
  DFFPOSX1 arr_reg_29__30_ ( .D(n7745), .CLK(clk), .Q(arr[987]) );
  DFFPOSX1 arr_reg_29__29_ ( .D(n7744), .CLK(clk), .Q(arr[986]) );
  DFFPOSX1 arr_reg_29__28_ ( .D(n7743), .CLK(clk), .Q(arr[985]) );
  DFFPOSX1 arr_reg_29__27_ ( .D(n7742), .CLK(clk), .Q(arr[984]) );
  DFFPOSX1 arr_reg_29__26_ ( .D(n7741), .CLK(clk), .Q(arr[983]) );
  DFFPOSX1 arr_reg_29__25_ ( .D(n7740), .CLK(clk), .Q(arr[982]) );
  DFFPOSX1 arr_reg_29__24_ ( .D(n7739), .CLK(clk), .Q(arr[981]) );
  DFFPOSX1 arr_reg_29__23_ ( .D(n7738), .CLK(clk), .Q(arr[980]) );
  DFFPOSX1 arr_reg_29__22_ ( .D(n7737), .CLK(clk), .Q(arr[979]) );
  DFFPOSX1 arr_reg_29__21_ ( .D(n7736), .CLK(clk), .Q(arr[978]) );
  DFFPOSX1 arr_reg_29__20_ ( .D(n7735), .CLK(clk), .Q(arr[977]) );
  DFFPOSX1 arr_reg_29__19_ ( .D(n7734), .CLK(clk), .Q(arr[976]) );
  DFFPOSX1 arr_reg_29__18_ ( .D(n7733), .CLK(clk), .Q(arr[975]) );
  DFFPOSX1 arr_reg_29__17_ ( .D(n7732), .CLK(clk), .Q(arr[974]) );
  DFFPOSX1 arr_reg_29__16_ ( .D(n7731), .CLK(clk), .Q(arr[973]) );
  DFFPOSX1 arr_reg_29__15_ ( .D(n7730), .CLK(clk), .Q(arr[972]) );
  DFFPOSX1 arr_reg_29__14_ ( .D(n7729), .CLK(clk), .Q(arr[971]) );
  DFFPOSX1 arr_reg_29__13_ ( .D(n7728), .CLK(clk), .Q(arr[970]) );
  DFFPOSX1 arr_reg_29__12_ ( .D(n7727), .CLK(clk), .Q(arr[969]) );
  DFFPOSX1 arr_reg_29__11_ ( .D(n7726), .CLK(clk), .Q(arr[968]) );
  DFFPOSX1 arr_reg_29__10_ ( .D(n7725), .CLK(clk), .Q(arr[967]) );
  DFFPOSX1 arr_reg_29__9_ ( .D(n7724), .CLK(clk), .Q(arr[966]) );
  DFFPOSX1 arr_reg_29__8_ ( .D(n7723), .CLK(clk), .Q(arr[965]) );
  DFFPOSX1 arr_reg_29__7_ ( .D(n7722), .CLK(clk), .Q(arr[964]) );
  DFFPOSX1 arr_reg_29__6_ ( .D(n7721), .CLK(clk), .Q(arr[963]) );
  DFFPOSX1 arr_reg_29__5_ ( .D(n7720), .CLK(clk), .Q(arr[962]) );
  DFFPOSX1 arr_reg_29__4_ ( .D(n7719), .CLK(clk), .Q(arr[961]) );
  DFFPOSX1 arr_reg_29__3_ ( .D(n7718), .CLK(clk), .Q(arr[960]) );
  DFFPOSX1 arr_reg_29__2_ ( .D(n7717), .CLK(clk), .Q(arr[959]) );
  DFFPOSX1 arr_reg_29__1_ ( .D(n7716), .CLK(clk), .Q(arr[958]) );
  DFFPOSX1 arr_reg_29__0_ ( .D(n7715), .CLK(clk), .Q(arr[957]) );
  DFFPOSX1 arr_reg_28__32_ ( .D(n7714), .CLK(clk), .Q(arr[956]) );
  DFFPOSX1 arr_reg_28__31_ ( .D(n7713), .CLK(clk), .Q(arr[955]) );
  DFFPOSX1 arr_reg_28__30_ ( .D(n7712), .CLK(clk), .Q(arr[954]) );
  DFFPOSX1 arr_reg_28__29_ ( .D(n7711), .CLK(clk), .Q(arr[953]) );
  DFFPOSX1 arr_reg_28__28_ ( .D(n7710), .CLK(clk), .Q(arr[952]) );
  DFFPOSX1 arr_reg_28__27_ ( .D(n7709), .CLK(clk), .Q(arr[951]) );
  DFFPOSX1 arr_reg_28__26_ ( .D(n7708), .CLK(clk), .Q(arr[950]) );
  DFFPOSX1 arr_reg_28__25_ ( .D(n7707), .CLK(clk), .Q(arr[949]) );
  DFFPOSX1 arr_reg_28__24_ ( .D(n7706), .CLK(clk), .Q(arr[948]) );
  DFFPOSX1 arr_reg_28__23_ ( .D(n7705), .CLK(clk), .Q(arr[947]) );
  DFFPOSX1 arr_reg_28__22_ ( .D(n7704), .CLK(clk), .Q(arr[946]) );
  DFFPOSX1 arr_reg_28__21_ ( .D(n7703), .CLK(clk), .Q(arr[945]) );
  DFFPOSX1 arr_reg_28__20_ ( .D(n7702), .CLK(clk), .Q(arr[944]) );
  DFFPOSX1 arr_reg_28__19_ ( .D(n7701), .CLK(clk), .Q(arr[943]) );
  DFFPOSX1 arr_reg_28__18_ ( .D(n7700), .CLK(clk), .Q(arr[942]) );
  DFFPOSX1 arr_reg_28__17_ ( .D(n7699), .CLK(clk), .Q(arr[941]) );
  DFFPOSX1 arr_reg_28__16_ ( .D(n7698), .CLK(clk), .Q(arr[940]) );
  DFFPOSX1 arr_reg_28__15_ ( .D(n7697), .CLK(clk), .Q(arr[939]) );
  DFFPOSX1 arr_reg_28__14_ ( .D(n7696), .CLK(clk), .Q(arr[938]) );
  DFFPOSX1 arr_reg_28__13_ ( .D(n7695), .CLK(clk), .Q(arr[937]) );
  DFFPOSX1 arr_reg_28__12_ ( .D(n7694), .CLK(clk), .Q(arr[936]) );
  DFFPOSX1 arr_reg_28__11_ ( .D(n7693), .CLK(clk), .Q(arr[935]) );
  DFFPOSX1 arr_reg_28__10_ ( .D(n7692), .CLK(clk), .Q(arr[934]) );
  DFFPOSX1 arr_reg_28__9_ ( .D(n7691), .CLK(clk), .Q(arr[933]) );
  DFFPOSX1 arr_reg_28__8_ ( .D(n7690), .CLK(clk), .Q(arr[932]) );
  DFFPOSX1 arr_reg_28__7_ ( .D(n7689), .CLK(clk), .Q(arr[931]) );
  DFFPOSX1 arr_reg_28__6_ ( .D(n7688), .CLK(clk), .Q(arr[930]) );
  DFFPOSX1 arr_reg_28__5_ ( .D(n7687), .CLK(clk), .Q(arr[929]) );
  DFFPOSX1 arr_reg_28__4_ ( .D(n7686), .CLK(clk), .Q(arr[928]) );
  DFFPOSX1 arr_reg_28__3_ ( .D(n7685), .CLK(clk), .Q(arr[927]) );
  DFFPOSX1 arr_reg_28__2_ ( .D(n7684), .CLK(clk), .Q(arr[926]) );
  DFFPOSX1 arr_reg_28__1_ ( .D(n7683), .CLK(clk), .Q(arr[925]) );
  DFFPOSX1 arr_reg_28__0_ ( .D(n7682), .CLK(clk), .Q(arr[924]) );
  DFFPOSX1 arr_reg_27__32_ ( .D(n7681), .CLK(clk), .Q(arr[923]) );
  DFFPOSX1 arr_reg_27__31_ ( .D(n7680), .CLK(clk), .Q(arr[922]) );
  DFFPOSX1 arr_reg_27__30_ ( .D(n7679), .CLK(clk), .Q(arr[921]) );
  DFFPOSX1 arr_reg_27__29_ ( .D(n7678), .CLK(clk), .Q(arr[920]) );
  DFFPOSX1 arr_reg_27__28_ ( .D(n7677), .CLK(clk), .Q(arr[919]) );
  DFFPOSX1 arr_reg_27__27_ ( .D(n7676), .CLK(clk), .Q(arr[918]) );
  DFFPOSX1 arr_reg_27__26_ ( .D(n7675), .CLK(clk), .Q(arr[917]) );
  DFFPOSX1 arr_reg_27__25_ ( .D(n7674), .CLK(clk), .Q(arr[916]) );
  DFFPOSX1 arr_reg_27__24_ ( .D(n7673), .CLK(clk), .Q(arr[915]) );
  DFFPOSX1 arr_reg_27__23_ ( .D(n7672), .CLK(clk), .Q(arr[914]) );
  DFFPOSX1 arr_reg_27__22_ ( .D(n7671), .CLK(clk), .Q(arr[913]) );
  DFFPOSX1 arr_reg_27__21_ ( .D(n7670), .CLK(clk), .Q(arr[912]) );
  DFFPOSX1 arr_reg_27__20_ ( .D(n7669), .CLK(clk), .Q(arr[911]) );
  DFFPOSX1 arr_reg_27__19_ ( .D(n7668), .CLK(clk), .Q(arr[910]) );
  DFFPOSX1 arr_reg_27__18_ ( .D(n7667), .CLK(clk), .Q(arr[909]) );
  DFFPOSX1 arr_reg_27__17_ ( .D(n7666), .CLK(clk), .Q(arr[908]) );
  DFFPOSX1 arr_reg_27__16_ ( .D(n7665), .CLK(clk), .Q(arr[907]) );
  DFFPOSX1 arr_reg_27__15_ ( .D(n7664), .CLK(clk), .Q(arr[906]) );
  DFFPOSX1 arr_reg_27__14_ ( .D(n7663), .CLK(clk), .Q(arr[905]) );
  DFFPOSX1 arr_reg_27__13_ ( .D(n7662), .CLK(clk), .Q(arr[904]) );
  DFFPOSX1 arr_reg_27__12_ ( .D(n7661), .CLK(clk), .Q(arr[903]) );
  DFFPOSX1 arr_reg_27__11_ ( .D(n7660), .CLK(clk), .Q(arr[902]) );
  DFFPOSX1 arr_reg_27__10_ ( .D(n7659), .CLK(clk), .Q(arr[901]) );
  DFFPOSX1 arr_reg_27__9_ ( .D(n7658), .CLK(clk), .Q(arr[900]) );
  DFFPOSX1 arr_reg_27__8_ ( .D(n7657), .CLK(clk), .Q(arr[899]) );
  DFFPOSX1 arr_reg_27__7_ ( .D(n7656), .CLK(clk), .Q(arr[898]) );
  DFFPOSX1 arr_reg_27__6_ ( .D(n7655), .CLK(clk), .Q(arr[897]) );
  DFFPOSX1 arr_reg_27__5_ ( .D(n7654), .CLK(clk), .Q(arr[896]) );
  DFFPOSX1 arr_reg_27__4_ ( .D(n7653), .CLK(clk), .Q(arr[895]) );
  DFFPOSX1 arr_reg_27__3_ ( .D(n7652), .CLK(clk), .Q(arr[894]) );
  DFFPOSX1 arr_reg_27__2_ ( .D(n7651), .CLK(clk), .Q(arr[893]) );
  DFFPOSX1 arr_reg_27__1_ ( .D(n7650), .CLK(clk), .Q(arr[892]) );
  DFFPOSX1 arr_reg_27__0_ ( .D(n7649), .CLK(clk), .Q(arr[891]) );
  DFFPOSX1 arr_reg_26__32_ ( .D(n7648), .CLK(clk), .Q(arr[890]) );
  DFFPOSX1 arr_reg_26__31_ ( .D(n7647), .CLK(clk), .Q(arr[889]) );
  DFFPOSX1 arr_reg_26__30_ ( .D(n7646), .CLK(clk), .Q(arr[888]) );
  DFFPOSX1 arr_reg_26__29_ ( .D(n7645), .CLK(clk), .Q(arr[887]) );
  DFFPOSX1 arr_reg_26__28_ ( .D(n7644), .CLK(clk), .Q(arr[886]) );
  DFFPOSX1 arr_reg_26__27_ ( .D(n7643), .CLK(clk), .Q(arr[885]) );
  DFFPOSX1 arr_reg_26__26_ ( .D(n7642), .CLK(clk), .Q(arr[884]) );
  DFFPOSX1 arr_reg_26__25_ ( .D(n7641), .CLK(clk), .Q(arr[883]) );
  DFFPOSX1 arr_reg_26__24_ ( .D(n7640), .CLK(clk), .Q(arr[882]) );
  DFFPOSX1 arr_reg_26__23_ ( .D(n7639), .CLK(clk), .Q(arr[881]) );
  DFFPOSX1 arr_reg_26__22_ ( .D(n7638), .CLK(clk), .Q(arr[880]) );
  DFFPOSX1 arr_reg_26__21_ ( .D(n7637), .CLK(clk), .Q(arr[879]) );
  DFFPOSX1 arr_reg_26__20_ ( .D(n7636), .CLK(clk), .Q(arr[878]) );
  DFFPOSX1 arr_reg_26__19_ ( .D(n7635), .CLK(clk), .Q(arr[877]) );
  DFFPOSX1 arr_reg_26__18_ ( .D(n7634), .CLK(clk), .Q(arr[876]) );
  DFFPOSX1 arr_reg_26__17_ ( .D(n7633), .CLK(clk), .Q(arr[875]) );
  DFFPOSX1 arr_reg_26__16_ ( .D(n7632), .CLK(clk), .Q(arr[874]) );
  DFFPOSX1 arr_reg_26__15_ ( .D(n7631), .CLK(clk), .Q(arr[873]) );
  DFFPOSX1 arr_reg_26__14_ ( .D(n7630), .CLK(clk), .Q(arr[872]) );
  DFFPOSX1 arr_reg_26__13_ ( .D(n7629), .CLK(clk), .Q(arr[871]) );
  DFFPOSX1 arr_reg_26__12_ ( .D(n7628), .CLK(clk), .Q(arr[870]) );
  DFFPOSX1 arr_reg_26__11_ ( .D(n7627), .CLK(clk), .Q(arr[869]) );
  DFFPOSX1 arr_reg_26__10_ ( .D(n7626), .CLK(clk), .Q(arr[868]) );
  DFFPOSX1 arr_reg_26__9_ ( .D(n7625), .CLK(clk), .Q(arr[867]) );
  DFFPOSX1 arr_reg_26__8_ ( .D(n7624), .CLK(clk), .Q(arr[866]) );
  DFFPOSX1 arr_reg_26__7_ ( .D(n7623), .CLK(clk), .Q(arr[865]) );
  DFFPOSX1 arr_reg_26__6_ ( .D(n7622), .CLK(clk), .Q(arr[864]) );
  DFFPOSX1 arr_reg_26__5_ ( .D(n7621), .CLK(clk), .Q(arr[863]) );
  DFFPOSX1 arr_reg_26__4_ ( .D(n7620), .CLK(clk), .Q(arr[862]) );
  DFFPOSX1 arr_reg_26__3_ ( .D(n7619), .CLK(clk), .Q(arr[861]) );
  DFFPOSX1 arr_reg_26__2_ ( .D(n7618), .CLK(clk), .Q(arr[860]) );
  DFFPOSX1 arr_reg_26__1_ ( .D(n7617), .CLK(clk), .Q(arr[859]) );
  DFFPOSX1 arr_reg_26__0_ ( .D(n7616), .CLK(clk), .Q(arr[858]) );
  DFFPOSX1 arr_reg_25__32_ ( .D(n7615), .CLK(clk), .Q(arr[857]) );
  DFFPOSX1 arr_reg_25__31_ ( .D(n7614), .CLK(clk), .Q(arr[856]) );
  DFFPOSX1 arr_reg_25__30_ ( .D(n7613), .CLK(clk), .Q(arr[855]) );
  DFFPOSX1 arr_reg_25__29_ ( .D(n7612), .CLK(clk), .Q(arr[854]) );
  DFFPOSX1 arr_reg_25__28_ ( .D(n7611), .CLK(clk), .Q(arr[853]) );
  DFFPOSX1 arr_reg_25__27_ ( .D(n7610), .CLK(clk), .Q(arr[852]) );
  DFFPOSX1 arr_reg_25__26_ ( .D(n7609), .CLK(clk), .Q(arr[851]) );
  DFFPOSX1 arr_reg_25__25_ ( .D(n7608), .CLK(clk), .Q(arr[850]) );
  DFFPOSX1 arr_reg_25__24_ ( .D(n7607), .CLK(clk), .Q(arr[849]) );
  DFFPOSX1 arr_reg_25__23_ ( .D(n7606), .CLK(clk), .Q(arr[848]) );
  DFFPOSX1 arr_reg_25__22_ ( .D(n7605), .CLK(clk), .Q(arr[847]) );
  DFFPOSX1 arr_reg_25__21_ ( .D(n7604), .CLK(clk), .Q(arr[846]) );
  DFFPOSX1 arr_reg_25__20_ ( .D(n7603), .CLK(clk), .Q(arr[845]) );
  DFFPOSX1 arr_reg_25__19_ ( .D(n7602), .CLK(clk), .Q(arr[844]) );
  DFFPOSX1 arr_reg_25__18_ ( .D(n7601), .CLK(clk), .Q(arr[843]) );
  DFFPOSX1 arr_reg_25__17_ ( .D(n7600), .CLK(clk), .Q(arr[842]) );
  DFFPOSX1 arr_reg_25__16_ ( .D(n7599), .CLK(clk), .Q(arr[841]) );
  DFFPOSX1 arr_reg_25__15_ ( .D(n7598), .CLK(clk), .Q(arr[840]) );
  DFFPOSX1 arr_reg_25__14_ ( .D(n7597), .CLK(clk), .Q(arr[839]) );
  DFFPOSX1 arr_reg_25__13_ ( .D(n7596), .CLK(clk), .Q(arr[838]) );
  DFFPOSX1 arr_reg_25__12_ ( .D(n7595), .CLK(clk), .Q(arr[837]) );
  DFFPOSX1 arr_reg_25__11_ ( .D(n7594), .CLK(clk), .Q(arr[836]) );
  DFFPOSX1 arr_reg_25__10_ ( .D(n7593), .CLK(clk), .Q(arr[835]) );
  DFFPOSX1 arr_reg_25__9_ ( .D(n7592), .CLK(clk), .Q(arr[834]) );
  DFFPOSX1 arr_reg_25__8_ ( .D(n7591), .CLK(clk), .Q(arr[833]) );
  DFFPOSX1 arr_reg_25__7_ ( .D(n7590), .CLK(clk), .Q(arr[832]) );
  DFFPOSX1 arr_reg_25__6_ ( .D(n7589), .CLK(clk), .Q(arr[831]) );
  DFFPOSX1 arr_reg_25__5_ ( .D(n7588), .CLK(clk), .Q(arr[830]) );
  DFFPOSX1 arr_reg_25__4_ ( .D(n7587), .CLK(clk), .Q(arr[829]) );
  DFFPOSX1 arr_reg_25__3_ ( .D(n7586), .CLK(clk), .Q(arr[828]) );
  DFFPOSX1 arr_reg_25__2_ ( .D(n7585), .CLK(clk), .Q(arr[827]) );
  DFFPOSX1 arr_reg_25__1_ ( .D(n7584), .CLK(clk), .Q(arr[826]) );
  DFFPOSX1 arr_reg_25__0_ ( .D(n7583), .CLK(clk), .Q(arr[825]) );
  DFFPOSX1 arr_reg_24__32_ ( .D(n7582), .CLK(clk), .Q(arr[824]) );
  DFFPOSX1 arr_reg_24__31_ ( .D(n7581), .CLK(clk), .Q(arr[823]) );
  DFFPOSX1 arr_reg_24__30_ ( .D(n7580), .CLK(clk), .Q(arr[822]) );
  DFFPOSX1 arr_reg_24__29_ ( .D(n7579), .CLK(clk), .Q(arr[821]) );
  DFFPOSX1 arr_reg_24__28_ ( .D(n7578), .CLK(clk), .Q(arr[820]) );
  DFFPOSX1 arr_reg_24__27_ ( .D(n7577), .CLK(clk), .Q(arr[819]) );
  DFFPOSX1 arr_reg_24__26_ ( .D(n7576), .CLK(clk), .Q(arr[818]) );
  DFFPOSX1 arr_reg_24__25_ ( .D(n7575), .CLK(clk), .Q(arr[817]) );
  DFFPOSX1 arr_reg_24__24_ ( .D(n7574), .CLK(clk), .Q(arr[816]) );
  DFFPOSX1 arr_reg_24__23_ ( .D(n7573), .CLK(clk), .Q(arr[815]) );
  DFFPOSX1 arr_reg_24__22_ ( .D(n7572), .CLK(clk), .Q(arr[814]) );
  DFFPOSX1 arr_reg_24__21_ ( .D(n7571), .CLK(clk), .Q(arr[813]) );
  DFFPOSX1 arr_reg_24__20_ ( .D(n7570), .CLK(clk), .Q(arr[812]) );
  DFFPOSX1 arr_reg_24__19_ ( .D(n7569), .CLK(clk), .Q(arr[811]) );
  DFFPOSX1 arr_reg_24__18_ ( .D(n7568), .CLK(clk), .Q(arr[810]) );
  DFFPOSX1 arr_reg_24__17_ ( .D(n7567), .CLK(clk), .Q(arr[809]) );
  DFFPOSX1 arr_reg_24__16_ ( .D(n7566), .CLK(clk), .Q(arr[808]) );
  DFFPOSX1 arr_reg_24__15_ ( .D(n7565), .CLK(clk), .Q(arr[807]) );
  DFFPOSX1 arr_reg_24__14_ ( .D(n7564), .CLK(clk), .Q(arr[806]) );
  DFFPOSX1 arr_reg_24__13_ ( .D(n7563), .CLK(clk), .Q(arr[805]) );
  DFFPOSX1 arr_reg_24__12_ ( .D(n7562), .CLK(clk), .Q(arr[804]) );
  DFFPOSX1 arr_reg_24__11_ ( .D(n7561), .CLK(clk), .Q(arr[803]) );
  DFFPOSX1 arr_reg_24__10_ ( .D(n7560), .CLK(clk), .Q(arr[802]) );
  DFFPOSX1 arr_reg_24__9_ ( .D(n7559), .CLK(clk), .Q(arr[801]) );
  DFFPOSX1 arr_reg_24__8_ ( .D(n7558), .CLK(clk), .Q(arr[800]) );
  DFFPOSX1 arr_reg_24__7_ ( .D(n7557), .CLK(clk), .Q(arr[799]) );
  DFFPOSX1 arr_reg_24__6_ ( .D(n7556), .CLK(clk), .Q(arr[798]) );
  DFFPOSX1 arr_reg_24__5_ ( .D(n7555), .CLK(clk), .Q(arr[797]) );
  DFFPOSX1 arr_reg_24__4_ ( .D(n7554), .CLK(clk), .Q(arr[796]) );
  DFFPOSX1 arr_reg_24__3_ ( .D(n7553), .CLK(clk), .Q(arr[795]) );
  DFFPOSX1 arr_reg_24__2_ ( .D(n7552), .CLK(clk), .Q(arr[794]) );
  DFFPOSX1 arr_reg_24__1_ ( .D(n7551), .CLK(clk), .Q(arr[793]) );
  DFFPOSX1 arr_reg_24__0_ ( .D(n7550), .CLK(clk), .Q(arr[792]) );
  DFFPOSX1 arr_reg_23__32_ ( .D(n7549), .CLK(clk), .Q(arr[791]) );
  DFFPOSX1 arr_reg_23__31_ ( .D(n7548), .CLK(clk), .Q(arr[790]) );
  DFFPOSX1 arr_reg_23__30_ ( .D(n7547), .CLK(clk), .Q(arr[789]) );
  DFFPOSX1 arr_reg_23__29_ ( .D(n7546), .CLK(clk), .Q(arr[788]) );
  DFFPOSX1 arr_reg_23__28_ ( .D(n7545), .CLK(clk), .Q(arr[787]) );
  DFFPOSX1 arr_reg_23__27_ ( .D(n7544), .CLK(clk), .Q(arr[786]) );
  DFFPOSX1 arr_reg_23__26_ ( .D(n7543), .CLK(clk), .Q(arr[785]) );
  DFFPOSX1 arr_reg_23__25_ ( .D(n7542), .CLK(clk), .Q(arr[784]) );
  DFFPOSX1 arr_reg_23__24_ ( .D(n7541), .CLK(clk), .Q(arr[783]) );
  DFFPOSX1 arr_reg_23__23_ ( .D(n7540), .CLK(clk), .Q(arr[782]) );
  DFFPOSX1 arr_reg_23__22_ ( .D(n7539), .CLK(clk), .Q(arr[781]) );
  DFFPOSX1 arr_reg_23__21_ ( .D(n7538), .CLK(clk), .Q(arr[780]) );
  DFFPOSX1 arr_reg_23__20_ ( .D(n7537), .CLK(clk), .Q(arr[779]) );
  DFFPOSX1 arr_reg_23__19_ ( .D(n7536), .CLK(clk), .Q(arr[778]) );
  DFFPOSX1 arr_reg_23__18_ ( .D(n7535), .CLK(clk), .Q(arr[777]) );
  DFFPOSX1 arr_reg_23__17_ ( .D(n7534), .CLK(clk), .Q(arr[776]) );
  DFFPOSX1 arr_reg_23__16_ ( .D(n7533), .CLK(clk), .Q(arr[775]) );
  DFFPOSX1 arr_reg_23__15_ ( .D(n7532), .CLK(clk), .Q(arr[774]) );
  DFFPOSX1 arr_reg_23__14_ ( .D(n7531), .CLK(clk), .Q(arr[773]) );
  DFFPOSX1 arr_reg_23__13_ ( .D(n7530), .CLK(clk), .Q(arr[772]) );
  DFFPOSX1 arr_reg_23__12_ ( .D(n7529), .CLK(clk), .Q(arr[771]) );
  DFFPOSX1 arr_reg_23__11_ ( .D(n7528), .CLK(clk), .Q(arr[770]) );
  DFFPOSX1 arr_reg_23__10_ ( .D(n7527), .CLK(clk), .Q(arr[769]) );
  DFFPOSX1 arr_reg_23__9_ ( .D(n7526), .CLK(clk), .Q(arr[768]) );
  DFFPOSX1 arr_reg_23__8_ ( .D(n7525), .CLK(clk), .Q(arr[767]) );
  DFFPOSX1 arr_reg_23__7_ ( .D(n7524), .CLK(clk), .Q(arr[766]) );
  DFFPOSX1 arr_reg_23__6_ ( .D(n7523), .CLK(clk), .Q(arr[765]) );
  DFFPOSX1 arr_reg_23__5_ ( .D(n7522), .CLK(clk), .Q(arr[764]) );
  DFFPOSX1 arr_reg_23__4_ ( .D(n7521), .CLK(clk), .Q(arr[763]) );
  DFFPOSX1 arr_reg_23__3_ ( .D(n7520), .CLK(clk), .Q(arr[762]) );
  DFFPOSX1 arr_reg_23__2_ ( .D(n7519), .CLK(clk), .Q(arr[761]) );
  DFFPOSX1 arr_reg_23__1_ ( .D(n7518), .CLK(clk), .Q(arr[760]) );
  DFFPOSX1 arr_reg_23__0_ ( .D(n7517), .CLK(clk), .Q(arr[759]) );
  DFFPOSX1 arr_reg_22__32_ ( .D(n7516), .CLK(clk), .Q(arr[758]) );
  DFFPOSX1 arr_reg_22__31_ ( .D(n7515), .CLK(clk), .Q(arr[757]) );
  DFFPOSX1 arr_reg_22__30_ ( .D(n7514), .CLK(clk), .Q(arr[756]) );
  DFFPOSX1 arr_reg_22__29_ ( .D(n7513), .CLK(clk), .Q(arr[755]) );
  DFFPOSX1 arr_reg_22__28_ ( .D(n7512), .CLK(clk), .Q(arr[754]) );
  DFFPOSX1 arr_reg_22__27_ ( .D(n7511), .CLK(clk), .Q(arr[753]) );
  DFFPOSX1 arr_reg_22__26_ ( .D(n7510), .CLK(clk), .Q(arr[752]) );
  DFFPOSX1 arr_reg_22__25_ ( .D(n7509), .CLK(clk), .Q(arr[751]) );
  DFFPOSX1 arr_reg_22__24_ ( .D(n7508), .CLK(clk), .Q(arr[750]) );
  DFFPOSX1 arr_reg_22__23_ ( .D(n7507), .CLK(clk), .Q(arr[749]) );
  DFFPOSX1 arr_reg_22__22_ ( .D(n7506), .CLK(clk), .Q(arr[748]) );
  DFFPOSX1 arr_reg_22__21_ ( .D(n7505), .CLK(clk), .Q(arr[747]) );
  DFFPOSX1 arr_reg_22__20_ ( .D(n7504), .CLK(clk), .Q(arr[746]) );
  DFFPOSX1 arr_reg_22__19_ ( .D(n7503), .CLK(clk), .Q(arr[745]) );
  DFFPOSX1 arr_reg_22__18_ ( .D(n7502), .CLK(clk), .Q(arr[744]) );
  DFFPOSX1 arr_reg_22__17_ ( .D(n7501), .CLK(clk), .Q(arr[743]) );
  DFFPOSX1 arr_reg_22__16_ ( .D(n7500), .CLK(clk), .Q(arr[742]) );
  DFFPOSX1 arr_reg_22__15_ ( .D(n7499), .CLK(clk), .Q(arr[741]) );
  DFFPOSX1 arr_reg_22__14_ ( .D(n7498), .CLK(clk), .Q(arr[740]) );
  DFFPOSX1 arr_reg_22__13_ ( .D(n7497), .CLK(clk), .Q(arr[739]) );
  DFFPOSX1 arr_reg_22__12_ ( .D(n7496), .CLK(clk), .Q(arr[738]) );
  DFFPOSX1 arr_reg_22__11_ ( .D(n7495), .CLK(clk), .Q(arr[737]) );
  DFFPOSX1 arr_reg_22__10_ ( .D(n7494), .CLK(clk), .Q(arr[736]) );
  DFFPOSX1 arr_reg_22__9_ ( .D(n7493), .CLK(clk), .Q(arr[735]) );
  DFFPOSX1 arr_reg_22__8_ ( .D(n7492), .CLK(clk), .Q(arr[734]) );
  DFFPOSX1 arr_reg_22__7_ ( .D(n7491), .CLK(clk), .Q(arr[733]) );
  DFFPOSX1 arr_reg_22__6_ ( .D(n7490), .CLK(clk), .Q(arr[732]) );
  DFFPOSX1 arr_reg_22__5_ ( .D(n7489), .CLK(clk), .Q(arr[731]) );
  DFFPOSX1 arr_reg_22__4_ ( .D(n7488), .CLK(clk), .Q(arr[730]) );
  DFFPOSX1 arr_reg_22__3_ ( .D(n7487), .CLK(clk), .Q(arr[729]) );
  DFFPOSX1 arr_reg_22__2_ ( .D(n7486), .CLK(clk), .Q(arr[728]) );
  DFFPOSX1 arr_reg_22__1_ ( .D(n7485), .CLK(clk), .Q(arr[727]) );
  DFFPOSX1 arr_reg_22__0_ ( .D(n7484), .CLK(clk), .Q(arr[726]) );
  DFFPOSX1 arr_reg_21__32_ ( .D(n7483), .CLK(clk), .Q(arr[725]) );
  DFFPOSX1 arr_reg_21__31_ ( .D(n7482), .CLK(clk), .Q(arr[724]) );
  DFFPOSX1 arr_reg_21__30_ ( .D(n7481), .CLK(clk), .Q(arr[723]) );
  DFFPOSX1 arr_reg_21__29_ ( .D(n7480), .CLK(clk), .Q(arr[722]) );
  DFFPOSX1 arr_reg_21__28_ ( .D(n7479), .CLK(clk), .Q(arr[721]) );
  DFFPOSX1 arr_reg_21__27_ ( .D(n7478), .CLK(clk), .Q(arr[720]) );
  DFFPOSX1 arr_reg_21__26_ ( .D(n7477), .CLK(clk), .Q(arr[719]) );
  DFFPOSX1 arr_reg_21__25_ ( .D(n7476), .CLK(clk), .Q(arr[718]) );
  DFFPOSX1 arr_reg_21__24_ ( .D(n7475), .CLK(clk), .Q(arr[717]) );
  DFFPOSX1 arr_reg_21__23_ ( .D(n7474), .CLK(clk), .Q(arr[716]) );
  DFFPOSX1 arr_reg_21__22_ ( .D(n7473), .CLK(clk), .Q(arr[715]) );
  DFFPOSX1 arr_reg_21__21_ ( .D(n7472), .CLK(clk), .Q(arr[714]) );
  DFFPOSX1 arr_reg_21__20_ ( .D(n7471), .CLK(clk), .Q(arr[713]) );
  DFFPOSX1 arr_reg_21__19_ ( .D(n7470), .CLK(clk), .Q(arr[712]) );
  DFFPOSX1 arr_reg_21__18_ ( .D(n7469), .CLK(clk), .Q(arr[711]) );
  DFFPOSX1 arr_reg_21__17_ ( .D(n7468), .CLK(clk), .Q(arr[710]) );
  DFFPOSX1 arr_reg_21__16_ ( .D(n7467), .CLK(clk), .Q(arr[709]) );
  DFFPOSX1 arr_reg_21__15_ ( .D(n7466), .CLK(clk), .Q(arr[708]) );
  DFFPOSX1 arr_reg_21__14_ ( .D(n7465), .CLK(clk), .Q(arr[707]) );
  DFFPOSX1 arr_reg_21__13_ ( .D(n7464), .CLK(clk), .Q(arr[706]) );
  DFFPOSX1 arr_reg_21__12_ ( .D(n7463), .CLK(clk), .Q(arr[705]) );
  DFFPOSX1 arr_reg_21__11_ ( .D(n7462), .CLK(clk), .Q(arr[704]) );
  DFFPOSX1 arr_reg_21__10_ ( .D(n7461), .CLK(clk), .Q(arr[703]) );
  DFFPOSX1 arr_reg_21__9_ ( .D(n7460), .CLK(clk), .Q(arr[702]) );
  DFFPOSX1 arr_reg_21__8_ ( .D(n7459), .CLK(clk), .Q(arr[701]) );
  DFFPOSX1 arr_reg_21__7_ ( .D(n7458), .CLK(clk), .Q(arr[700]) );
  DFFPOSX1 arr_reg_21__6_ ( .D(n7457), .CLK(clk), .Q(arr[699]) );
  DFFPOSX1 arr_reg_21__5_ ( .D(n7456), .CLK(clk), .Q(arr[698]) );
  DFFPOSX1 arr_reg_21__4_ ( .D(n7455), .CLK(clk), .Q(arr[697]) );
  DFFPOSX1 arr_reg_21__3_ ( .D(n7454), .CLK(clk), .Q(arr[696]) );
  DFFPOSX1 arr_reg_21__2_ ( .D(n7453), .CLK(clk), .Q(arr[695]) );
  DFFPOSX1 arr_reg_21__1_ ( .D(n7452), .CLK(clk), .Q(arr[694]) );
  DFFPOSX1 arr_reg_21__0_ ( .D(n7451), .CLK(clk), .Q(arr[693]) );
  DFFPOSX1 arr_reg_20__32_ ( .D(n7450), .CLK(clk), .Q(arr[692]) );
  DFFPOSX1 arr_reg_20__31_ ( .D(n7449), .CLK(clk), .Q(arr[691]) );
  DFFPOSX1 arr_reg_20__30_ ( .D(n7448), .CLK(clk), .Q(arr[690]) );
  DFFPOSX1 arr_reg_20__29_ ( .D(n7447), .CLK(clk), .Q(arr[689]) );
  DFFPOSX1 arr_reg_20__28_ ( .D(n7446), .CLK(clk), .Q(arr[688]) );
  DFFPOSX1 arr_reg_20__27_ ( .D(n7445), .CLK(clk), .Q(arr[687]) );
  DFFPOSX1 arr_reg_20__26_ ( .D(n7444), .CLK(clk), .Q(arr[686]) );
  DFFPOSX1 arr_reg_20__25_ ( .D(n7443), .CLK(clk), .Q(arr[685]) );
  DFFPOSX1 arr_reg_20__24_ ( .D(n7442), .CLK(clk), .Q(arr[684]) );
  DFFPOSX1 arr_reg_20__23_ ( .D(n7441), .CLK(clk), .Q(arr[683]) );
  DFFPOSX1 arr_reg_20__22_ ( .D(n7440), .CLK(clk), .Q(arr[682]) );
  DFFPOSX1 arr_reg_20__21_ ( .D(n7439), .CLK(clk), .Q(arr[681]) );
  DFFPOSX1 arr_reg_20__20_ ( .D(n7438), .CLK(clk), .Q(arr[680]) );
  DFFPOSX1 arr_reg_20__19_ ( .D(n7437), .CLK(clk), .Q(arr[679]) );
  DFFPOSX1 arr_reg_20__18_ ( .D(n7436), .CLK(clk), .Q(arr[678]) );
  DFFPOSX1 arr_reg_20__17_ ( .D(n7435), .CLK(clk), .Q(arr[677]) );
  DFFPOSX1 arr_reg_20__16_ ( .D(n7434), .CLK(clk), .Q(arr[676]) );
  DFFPOSX1 arr_reg_20__15_ ( .D(n7433), .CLK(clk), .Q(arr[675]) );
  DFFPOSX1 arr_reg_20__14_ ( .D(n7432), .CLK(clk), .Q(arr[674]) );
  DFFPOSX1 arr_reg_20__13_ ( .D(n7431), .CLK(clk), .Q(arr[673]) );
  DFFPOSX1 arr_reg_20__12_ ( .D(n7430), .CLK(clk), .Q(arr[672]) );
  DFFPOSX1 arr_reg_20__11_ ( .D(n7429), .CLK(clk), .Q(arr[671]) );
  DFFPOSX1 arr_reg_20__10_ ( .D(n7428), .CLK(clk), .Q(arr[670]) );
  DFFPOSX1 arr_reg_20__9_ ( .D(n7427), .CLK(clk), .Q(arr[669]) );
  DFFPOSX1 arr_reg_20__8_ ( .D(n7426), .CLK(clk), .Q(arr[668]) );
  DFFPOSX1 arr_reg_20__7_ ( .D(n7425), .CLK(clk), .Q(arr[667]) );
  DFFPOSX1 arr_reg_20__6_ ( .D(n7424), .CLK(clk), .Q(arr[666]) );
  DFFPOSX1 arr_reg_20__5_ ( .D(n7423), .CLK(clk), .Q(arr[665]) );
  DFFPOSX1 arr_reg_20__4_ ( .D(n7422), .CLK(clk), .Q(arr[664]) );
  DFFPOSX1 arr_reg_20__3_ ( .D(n7421), .CLK(clk), .Q(arr[663]) );
  DFFPOSX1 arr_reg_20__2_ ( .D(n7420), .CLK(clk), .Q(arr[662]) );
  DFFPOSX1 arr_reg_20__1_ ( .D(n7419), .CLK(clk), .Q(arr[661]) );
  DFFPOSX1 arr_reg_20__0_ ( .D(n7418), .CLK(clk), .Q(arr[660]) );
  DFFPOSX1 arr_reg_19__32_ ( .D(n7417), .CLK(clk), .Q(arr[659]) );
  DFFPOSX1 arr_reg_19__31_ ( .D(n7416), .CLK(clk), .Q(arr[658]) );
  DFFPOSX1 arr_reg_19__30_ ( .D(n7415), .CLK(clk), .Q(arr[657]) );
  DFFPOSX1 arr_reg_19__29_ ( .D(n7414), .CLK(clk), .Q(arr[656]) );
  DFFPOSX1 arr_reg_19__28_ ( .D(n7413), .CLK(clk), .Q(arr[655]) );
  DFFPOSX1 arr_reg_19__27_ ( .D(n7412), .CLK(clk), .Q(arr[654]) );
  DFFPOSX1 arr_reg_19__26_ ( .D(n7411), .CLK(clk), .Q(arr[653]) );
  DFFPOSX1 arr_reg_19__25_ ( .D(n7410), .CLK(clk), .Q(arr[652]) );
  DFFPOSX1 arr_reg_19__24_ ( .D(n7409), .CLK(clk), .Q(arr[651]) );
  DFFPOSX1 arr_reg_19__23_ ( .D(n7408), .CLK(clk), .Q(arr[650]) );
  DFFPOSX1 arr_reg_19__22_ ( .D(n7407), .CLK(clk), .Q(arr[649]) );
  DFFPOSX1 arr_reg_19__21_ ( .D(n7406), .CLK(clk), .Q(arr[648]) );
  DFFPOSX1 arr_reg_19__20_ ( .D(n7405), .CLK(clk), .Q(arr[647]) );
  DFFPOSX1 arr_reg_19__19_ ( .D(n7404), .CLK(clk), .Q(arr[646]) );
  DFFPOSX1 arr_reg_19__18_ ( .D(n7403), .CLK(clk), .Q(arr[645]) );
  DFFPOSX1 arr_reg_19__17_ ( .D(n7402), .CLK(clk), .Q(arr[644]) );
  DFFPOSX1 arr_reg_19__16_ ( .D(n7401), .CLK(clk), .Q(arr[643]) );
  DFFPOSX1 arr_reg_19__15_ ( .D(n7400), .CLK(clk), .Q(arr[642]) );
  DFFPOSX1 arr_reg_19__14_ ( .D(n7399), .CLK(clk), .Q(arr[641]) );
  DFFPOSX1 arr_reg_19__13_ ( .D(n7398), .CLK(clk), .Q(arr[640]) );
  DFFPOSX1 arr_reg_19__12_ ( .D(n7397), .CLK(clk), .Q(arr[639]) );
  DFFPOSX1 arr_reg_19__11_ ( .D(n7396), .CLK(clk), .Q(arr[638]) );
  DFFPOSX1 arr_reg_19__10_ ( .D(n7395), .CLK(clk), .Q(arr[637]) );
  DFFPOSX1 arr_reg_19__9_ ( .D(n7394), .CLK(clk), .Q(arr[636]) );
  DFFPOSX1 arr_reg_19__8_ ( .D(n7393), .CLK(clk), .Q(arr[635]) );
  DFFPOSX1 arr_reg_19__7_ ( .D(n7392), .CLK(clk), .Q(arr[634]) );
  DFFPOSX1 arr_reg_19__6_ ( .D(n7391), .CLK(clk), .Q(arr[633]) );
  DFFPOSX1 arr_reg_19__5_ ( .D(n7390), .CLK(clk), .Q(arr[632]) );
  DFFPOSX1 arr_reg_19__4_ ( .D(n7389), .CLK(clk), .Q(arr[631]) );
  DFFPOSX1 arr_reg_19__3_ ( .D(n7388), .CLK(clk), .Q(arr[630]) );
  DFFPOSX1 arr_reg_19__2_ ( .D(n7387), .CLK(clk), .Q(arr[629]) );
  DFFPOSX1 arr_reg_19__1_ ( .D(n7386), .CLK(clk), .Q(arr[628]) );
  DFFPOSX1 arr_reg_19__0_ ( .D(n7385), .CLK(clk), .Q(arr[627]) );
  DFFPOSX1 arr_reg_18__32_ ( .D(n7384), .CLK(clk), .Q(arr[626]) );
  DFFPOSX1 arr_reg_18__31_ ( .D(n7383), .CLK(clk), .Q(arr[625]) );
  DFFPOSX1 arr_reg_18__30_ ( .D(n7382), .CLK(clk), .Q(arr[624]) );
  DFFPOSX1 arr_reg_18__29_ ( .D(n7381), .CLK(clk), .Q(arr[623]) );
  DFFPOSX1 arr_reg_18__28_ ( .D(n7380), .CLK(clk), .Q(arr[622]) );
  DFFPOSX1 arr_reg_18__27_ ( .D(n7379), .CLK(clk), .Q(arr[621]) );
  DFFPOSX1 arr_reg_18__26_ ( .D(n7378), .CLK(clk), .Q(arr[620]) );
  DFFPOSX1 arr_reg_18__25_ ( .D(n7377), .CLK(clk), .Q(arr[619]) );
  DFFPOSX1 arr_reg_18__24_ ( .D(n7376), .CLK(clk), .Q(arr[618]) );
  DFFPOSX1 arr_reg_18__23_ ( .D(n7375), .CLK(clk), .Q(arr[617]) );
  DFFPOSX1 arr_reg_18__22_ ( .D(n7374), .CLK(clk), .Q(arr[616]) );
  DFFPOSX1 arr_reg_18__21_ ( .D(n7373), .CLK(clk), .Q(arr[615]) );
  DFFPOSX1 arr_reg_18__20_ ( .D(n7372), .CLK(clk), .Q(arr[614]) );
  DFFPOSX1 arr_reg_18__19_ ( .D(n7371), .CLK(clk), .Q(arr[613]) );
  DFFPOSX1 arr_reg_18__18_ ( .D(n7370), .CLK(clk), .Q(arr[612]) );
  DFFPOSX1 arr_reg_18__17_ ( .D(n7369), .CLK(clk), .Q(arr[611]) );
  DFFPOSX1 arr_reg_18__16_ ( .D(n7368), .CLK(clk), .Q(arr[610]) );
  DFFPOSX1 arr_reg_18__15_ ( .D(n7367), .CLK(clk), .Q(arr[609]) );
  DFFPOSX1 arr_reg_18__14_ ( .D(n7366), .CLK(clk), .Q(arr[608]) );
  DFFPOSX1 arr_reg_18__13_ ( .D(n7365), .CLK(clk), .Q(arr[607]) );
  DFFPOSX1 arr_reg_18__12_ ( .D(n7364), .CLK(clk), .Q(arr[606]) );
  DFFPOSX1 arr_reg_18__11_ ( .D(n7363), .CLK(clk), .Q(arr[605]) );
  DFFPOSX1 arr_reg_18__10_ ( .D(n7362), .CLK(clk), .Q(arr[604]) );
  DFFPOSX1 arr_reg_18__9_ ( .D(n7361), .CLK(clk), .Q(arr[603]) );
  DFFPOSX1 arr_reg_18__8_ ( .D(n7360), .CLK(clk), .Q(arr[602]) );
  DFFPOSX1 arr_reg_18__7_ ( .D(n7359), .CLK(clk), .Q(arr[601]) );
  DFFPOSX1 arr_reg_18__6_ ( .D(n7358), .CLK(clk), .Q(arr[600]) );
  DFFPOSX1 arr_reg_18__5_ ( .D(n7357), .CLK(clk), .Q(arr[599]) );
  DFFPOSX1 arr_reg_18__4_ ( .D(n7356), .CLK(clk), .Q(arr[598]) );
  DFFPOSX1 arr_reg_18__3_ ( .D(n7355), .CLK(clk), .Q(arr[597]) );
  DFFPOSX1 arr_reg_18__2_ ( .D(n7354), .CLK(clk), .Q(arr[596]) );
  DFFPOSX1 arr_reg_18__1_ ( .D(n7353), .CLK(clk), .Q(arr[595]) );
  DFFPOSX1 arr_reg_18__0_ ( .D(n7352), .CLK(clk), .Q(arr[594]) );
  DFFPOSX1 arr_reg_17__32_ ( .D(n7351), .CLK(clk), .Q(arr[593]) );
  DFFPOSX1 arr_reg_17__31_ ( .D(n7350), .CLK(clk), .Q(arr[592]) );
  DFFPOSX1 arr_reg_17__30_ ( .D(n7349), .CLK(clk), .Q(arr[591]) );
  DFFPOSX1 arr_reg_17__29_ ( .D(n7348), .CLK(clk), .Q(arr[590]) );
  DFFPOSX1 arr_reg_17__28_ ( .D(n7347), .CLK(clk), .Q(arr[589]) );
  DFFPOSX1 arr_reg_17__27_ ( .D(n7346), .CLK(clk), .Q(arr[588]) );
  DFFPOSX1 arr_reg_17__26_ ( .D(n7345), .CLK(clk), .Q(arr[587]) );
  DFFPOSX1 arr_reg_17__25_ ( .D(n7344), .CLK(clk), .Q(arr[586]) );
  DFFPOSX1 arr_reg_17__24_ ( .D(n7343), .CLK(clk), .Q(arr[585]) );
  DFFPOSX1 arr_reg_17__23_ ( .D(n7342), .CLK(clk), .Q(arr[584]) );
  DFFPOSX1 arr_reg_17__22_ ( .D(n7341), .CLK(clk), .Q(arr[583]) );
  DFFPOSX1 arr_reg_17__21_ ( .D(n7340), .CLK(clk), .Q(arr[582]) );
  DFFPOSX1 arr_reg_17__20_ ( .D(n7339), .CLK(clk), .Q(arr[581]) );
  DFFPOSX1 arr_reg_17__19_ ( .D(n7338), .CLK(clk), .Q(arr[580]) );
  DFFPOSX1 arr_reg_17__18_ ( .D(n7337), .CLK(clk), .Q(arr[579]) );
  DFFPOSX1 arr_reg_17__17_ ( .D(n7336), .CLK(clk), .Q(arr[578]) );
  DFFPOSX1 arr_reg_17__16_ ( .D(n7335), .CLK(clk), .Q(arr[577]) );
  DFFPOSX1 arr_reg_17__15_ ( .D(n7334), .CLK(clk), .Q(arr[576]) );
  DFFPOSX1 arr_reg_17__14_ ( .D(n7333), .CLK(clk), .Q(arr[575]) );
  DFFPOSX1 arr_reg_17__13_ ( .D(n7332), .CLK(clk), .Q(arr[574]) );
  DFFPOSX1 arr_reg_17__12_ ( .D(n7331), .CLK(clk), .Q(arr[573]) );
  DFFPOSX1 arr_reg_17__11_ ( .D(n7330), .CLK(clk), .Q(arr[572]) );
  DFFPOSX1 arr_reg_17__10_ ( .D(n7329), .CLK(clk), .Q(arr[571]) );
  DFFPOSX1 arr_reg_17__9_ ( .D(n7328), .CLK(clk), .Q(arr[570]) );
  DFFPOSX1 arr_reg_17__8_ ( .D(n7327), .CLK(clk), .Q(arr[569]) );
  DFFPOSX1 arr_reg_17__7_ ( .D(n7326), .CLK(clk), .Q(arr[568]) );
  DFFPOSX1 arr_reg_17__6_ ( .D(n7325), .CLK(clk), .Q(arr[567]) );
  DFFPOSX1 arr_reg_17__5_ ( .D(n7324), .CLK(clk), .Q(arr[566]) );
  DFFPOSX1 arr_reg_17__4_ ( .D(n7323), .CLK(clk), .Q(arr[565]) );
  DFFPOSX1 arr_reg_17__3_ ( .D(n7322), .CLK(clk), .Q(arr[564]) );
  DFFPOSX1 arr_reg_17__2_ ( .D(n7321), .CLK(clk), .Q(arr[563]) );
  DFFPOSX1 arr_reg_17__1_ ( .D(n7320), .CLK(clk), .Q(arr[562]) );
  DFFPOSX1 arr_reg_17__0_ ( .D(n7319), .CLK(clk), .Q(arr[561]) );
  DFFPOSX1 arr_reg_16__32_ ( .D(n7318), .CLK(clk), .Q(arr[560]) );
  DFFPOSX1 arr_reg_16__31_ ( .D(n7317), .CLK(clk), .Q(arr[559]) );
  DFFPOSX1 arr_reg_16__30_ ( .D(n7316), .CLK(clk), .Q(arr[558]) );
  DFFPOSX1 arr_reg_16__29_ ( .D(n7315), .CLK(clk), .Q(arr[557]) );
  DFFPOSX1 arr_reg_16__28_ ( .D(n7314), .CLK(clk), .Q(arr[556]) );
  DFFPOSX1 arr_reg_16__27_ ( .D(n7313), .CLK(clk), .Q(arr[555]) );
  DFFPOSX1 arr_reg_16__26_ ( .D(n7312), .CLK(clk), .Q(arr[554]) );
  DFFPOSX1 arr_reg_16__25_ ( .D(n7311), .CLK(clk), .Q(arr[553]) );
  DFFPOSX1 arr_reg_16__24_ ( .D(n7310), .CLK(clk), .Q(arr[552]) );
  DFFPOSX1 arr_reg_16__23_ ( .D(n7309), .CLK(clk), .Q(arr[551]) );
  DFFPOSX1 arr_reg_16__22_ ( .D(n7308), .CLK(clk), .Q(arr[550]) );
  DFFPOSX1 arr_reg_16__21_ ( .D(n7307), .CLK(clk), .Q(arr[549]) );
  DFFPOSX1 arr_reg_16__20_ ( .D(n7306), .CLK(clk), .Q(arr[548]) );
  DFFPOSX1 arr_reg_16__19_ ( .D(n7305), .CLK(clk), .Q(arr[547]) );
  DFFPOSX1 arr_reg_16__18_ ( .D(n7304), .CLK(clk), .Q(arr[546]) );
  DFFPOSX1 arr_reg_16__17_ ( .D(n7303), .CLK(clk), .Q(arr[545]) );
  DFFPOSX1 arr_reg_16__16_ ( .D(n7302), .CLK(clk), .Q(arr[544]) );
  DFFPOSX1 arr_reg_16__15_ ( .D(n7301), .CLK(clk), .Q(arr[543]) );
  DFFPOSX1 arr_reg_16__14_ ( .D(n7300), .CLK(clk), .Q(arr[542]) );
  DFFPOSX1 arr_reg_16__13_ ( .D(n7299), .CLK(clk), .Q(arr[541]) );
  DFFPOSX1 arr_reg_16__12_ ( .D(n7298), .CLK(clk), .Q(arr[540]) );
  DFFPOSX1 arr_reg_16__11_ ( .D(n7297), .CLK(clk), .Q(arr[539]) );
  DFFPOSX1 arr_reg_16__10_ ( .D(n7296), .CLK(clk), .Q(arr[538]) );
  DFFPOSX1 arr_reg_16__9_ ( .D(n7295), .CLK(clk), .Q(arr[537]) );
  DFFPOSX1 arr_reg_16__8_ ( .D(n7294), .CLK(clk), .Q(arr[536]) );
  DFFPOSX1 arr_reg_16__7_ ( .D(n7293), .CLK(clk), .Q(arr[535]) );
  DFFPOSX1 arr_reg_16__6_ ( .D(n7292), .CLK(clk), .Q(arr[534]) );
  DFFPOSX1 arr_reg_16__5_ ( .D(n7291), .CLK(clk), .Q(arr[533]) );
  DFFPOSX1 arr_reg_16__4_ ( .D(n7290), .CLK(clk), .Q(arr[532]) );
  DFFPOSX1 arr_reg_16__3_ ( .D(n7289), .CLK(clk), .Q(arr[531]) );
  DFFPOSX1 arr_reg_16__2_ ( .D(n7288), .CLK(clk), .Q(arr[530]) );
  DFFPOSX1 arr_reg_16__1_ ( .D(n7287), .CLK(clk), .Q(arr[529]) );
  DFFPOSX1 arr_reg_16__0_ ( .D(n7286), .CLK(clk), .Q(arr[528]) );
  DFFPOSX1 arr_reg_15__32_ ( .D(n7285), .CLK(clk), .Q(arr[527]) );
  DFFPOSX1 arr_reg_15__31_ ( .D(n7284), .CLK(clk), .Q(arr[526]) );
  DFFPOSX1 arr_reg_15__30_ ( .D(n7283), .CLK(clk), .Q(arr[525]) );
  DFFPOSX1 arr_reg_15__29_ ( .D(n7282), .CLK(clk), .Q(arr[524]) );
  DFFPOSX1 arr_reg_15__28_ ( .D(n7281), .CLK(clk), .Q(arr[523]) );
  DFFPOSX1 arr_reg_15__27_ ( .D(n7280), .CLK(clk), .Q(arr[522]) );
  DFFPOSX1 arr_reg_15__26_ ( .D(n7279), .CLK(clk), .Q(arr[521]) );
  DFFPOSX1 arr_reg_15__25_ ( .D(n7278), .CLK(clk), .Q(arr[520]) );
  DFFPOSX1 arr_reg_15__24_ ( .D(n7277), .CLK(clk), .Q(arr[519]) );
  DFFPOSX1 arr_reg_15__23_ ( .D(n7276), .CLK(clk), .Q(arr[518]) );
  DFFPOSX1 arr_reg_15__22_ ( .D(n7275), .CLK(clk), .Q(arr[517]) );
  DFFPOSX1 arr_reg_15__21_ ( .D(n7274), .CLK(clk), .Q(arr[516]) );
  DFFPOSX1 arr_reg_15__20_ ( .D(n7273), .CLK(clk), .Q(arr[515]) );
  DFFPOSX1 arr_reg_15__19_ ( .D(n7272), .CLK(clk), .Q(arr[514]) );
  DFFPOSX1 arr_reg_15__18_ ( .D(n7271), .CLK(clk), .Q(arr[513]) );
  DFFPOSX1 arr_reg_15__17_ ( .D(n7270), .CLK(clk), .Q(arr[512]) );
  DFFPOSX1 arr_reg_15__16_ ( .D(n7269), .CLK(clk), .Q(arr[511]) );
  DFFPOSX1 arr_reg_15__15_ ( .D(n7268), .CLK(clk), .Q(arr[510]) );
  DFFPOSX1 arr_reg_15__14_ ( .D(n7267), .CLK(clk), .Q(arr[509]) );
  DFFPOSX1 arr_reg_15__13_ ( .D(n7266), .CLK(clk), .Q(arr[508]) );
  DFFPOSX1 arr_reg_15__12_ ( .D(n7265), .CLK(clk), .Q(arr[507]) );
  DFFPOSX1 arr_reg_15__11_ ( .D(n7264), .CLK(clk), .Q(arr[506]) );
  DFFPOSX1 arr_reg_15__10_ ( .D(n7263), .CLK(clk), .Q(arr[505]) );
  DFFPOSX1 arr_reg_15__9_ ( .D(n7262), .CLK(clk), .Q(arr[504]) );
  DFFPOSX1 arr_reg_15__8_ ( .D(n7261), .CLK(clk), .Q(arr[503]) );
  DFFPOSX1 arr_reg_15__7_ ( .D(n7260), .CLK(clk), .Q(arr[502]) );
  DFFPOSX1 arr_reg_15__6_ ( .D(n7259), .CLK(clk), .Q(arr[501]) );
  DFFPOSX1 arr_reg_15__5_ ( .D(n7258), .CLK(clk), .Q(arr[500]) );
  DFFPOSX1 arr_reg_15__4_ ( .D(n7257), .CLK(clk), .Q(arr[499]) );
  DFFPOSX1 arr_reg_15__3_ ( .D(n7256), .CLK(clk), .Q(arr[498]) );
  DFFPOSX1 arr_reg_15__2_ ( .D(n7255), .CLK(clk), .Q(arr[497]) );
  DFFPOSX1 arr_reg_15__1_ ( .D(n7254), .CLK(clk), .Q(arr[496]) );
  DFFPOSX1 arr_reg_15__0_ ( .D(n7253), .CLK(clk), .Q(arr[495]) );
  DFFPOSX1 arr_reg_14__32_ ( .D(n7252), .CLK(clk), .Q(arr[494]) );
  DFFPOSX1 arr_reg_14__31_ ( .D(n7251), .CLK(clk), .Q(arr[493]) );
  DFFPOSX1 arr_reg_14__30_ ( .D(n7250), .CLK(clk), .Q(arr[492]) );
  DFFPOSX1 arr_reg_14__29_ ( .D(n7249), .CLK(clk), .Q(arr[491]) );
  DFFPOSX1 arr_reg_14__28_ ( .D(n7248), .CLK(clk), .Q(arr[490]) );
  DFFPOSX1 arr_reg_14__27_ ( .D(n7247), .CLK(clk), .Q(arr[489]) );
  DFFPOSX1 arr_reg_14__26_ ( .D(n7246), .CLK(clk), .Q(arr[488]) );
  DFFPOSX1 arr_reg_14__25_ ( .D(n7245), .CLK(clk), .Q(arr[487]) );
  DFFPOSX1 arr_reg_14__24_ ( .D(n7244), .CLK(clk), .Q(arr[486]) );
  DFFPOSX1 arr_reg_14__23_ ( .D(n7243), .CLK(clk), .Q(arr[485]) );
  DFFPOSX1 arr_reg_14__22_ ( .D(n7242), .CLK(clk), .Q(arr[484]) );
  DFFPOSX1 arr_reg_14__21_ ( .D(n7241), .CLK(clk), .Q(arr[483]) );
  DFFPOSX1 arr_reg_14__20_ ( .D(n7240), .CLK(clk), .Q(arr[482]) );
  DFFPOSX1 arr_reg_14__19_ ( .D(n7239), .CLK(clk), .Q(arr[481]) );
  DFFPOSX1 arr_reg_14__18_ ( .D(n7238), .CLK(clk), .Q(arr[480]) );
  DFFPOSX1 arr_reg_14__17_ ( .D(n7237), .CLK(clk), .Q(arr[479]) );
  DFFPOSX1 arr_reg_14__16_ ( .D(n7236), .CLK(clk), .Q(arr[478]) );
  DFFPOSX1 arr_reg_14__15_ ( .D(n7235), .CLK(clk), .Q(arr[477]) );
  DFFPOSX1 arr_reg_14__14_ ( .D(n7234), .CLK(clk), .Q(arr[476]) );
  DFFPOSX1 arr_reg_14__13_ ( .D(n7233), .CLK(clk), .Q(arr[475]) );
  DFFPOSX1 arr_reg_14__12_ ( .D(n7232), .CLK(clk), .Q(arr[474]) );
  DFFPOSX1 arr_reg_14__11_ ( .D(n7231), .CLK(clk), .Q(arr[473]) );
  DFFPOSX1 arr_reg_14__10_ ( .D(n7230), .CLK(clk), .Q(arr[472]) );
  DFFPOSX1 arr_reg_14__9_ ( .D(n7229), .CLK(clk), .Q(arr[471]) );
  DFFPOSX1 arr_reg_14__8_ ( .D(n7228), .CLK(clk), .Q(arr[470]) );
  DFFPOSX1 arr_reg_14__7_ ( .D(n7227), .CLK(clk), .Q(arr[469]) );
  DFFPOSX1 arr_reg_14__6_ ( .D(n7226), .CLK(clk), .Q(arr[468]) );
  DFFPOSX1 arr_reg_14__5_ ( .D(n7225), .CLK(clk), .Q(arr[467]) );
  DFFPOSX1 arr_reg_14__4_ ( .D(n7224), .CLK(clk), .Q(arr[466]) );
  DFFPOSX1 arr_reg_14__3_ ( .D(n7223), .CLK(clk), .Q(arr[465]) );
  DFFPOSX1 arr_reg_14__2_ ( .D(n7222), .CLK(clk), .Q(arr[464]) );
  DFFPOSX1 arr_reg_14__1_ ( .D(n7221), .CLK(clk), .Q(arr[463]) );
  DFFPOSX1 arr_reg_14__0_ ( .D(n7220), .CLK(clk), .Q(arr[462]) );
  DFFPOSX1 arr_reg_13__32_ ( .D(n7219), .CLK(clk), .Q(arr[461]) );
  DFFPOSX1 arr_reg_13__31_ ( .D(n7218), .CLK(clk), .Q(arr[460]) );
  DFFPOSX1 arr_reg_13__30_ ( .D(n7217), .CLK(clk), .Q(arr[459]) );
  DFFPOSX1 arr_reg_13__29_ ( .D(n7216), .CLK(clk), .Q(arr[458]) );
  DFFPOSX1 arr_reg_13__28_ ( .D(n7215), .CLK(clk), .Q(arr[457]) );
  DFFPOSX1 arr_reg_13__27_ ( .D(n7214), .CLK(clk), .Q(arr[456]) );
  DFFPOSX1 arr_reg_13__26_ ( .D(n7213), .CLK(clk), .Q(arr[455]) );
  DFFPOSX1 arr_reg_13__25_ ( .D(n7212), .CLK(clk), .Q(arr[454]) );
  DFFPOSX1 arr_reg_13__24_ ( .D(n7211), .CLK(clk), .Q(arr[453]) );
  DFFPOSX1 arr_reg_13__23_ ( .D(n7210), .CLK(clk), .Q(arr[452]) );
  DFFPOSX1 arr_reg_13__22_ ( .D(n7209), .CLK(clk), .Q(arr[451]) );
  DFFPOSX1 arr_reg_13__21_ ( .D(n7208), .CLK(clk), .Q(arr[450]) );
  DFFPOSX1 arr_reg_13__20_ ( .D(n7207), .CLK(clk), .Q(arr[449]) );
  DFFPOSX1 arr_reg_13__19_ ( .D(n7206), .CLK(clk), .Q(arr[448]) );
  DFFPOSX1 arr_reg_13__18_ ( .D(n7205), .CLK(clk), .Q(arr[447]) );
  DFFPOSX1 arr_reg_13__17_ ( .D(n7204), .CLK(clk), .Q(arr[446]) );
  DFFPOSX1 arr_reg_13__16_ ( .D(n7203), .CLK(clk), .Q(arr[445]) );
  DFFPOSX1 arr_reg_13__15_ ( .D(n7202), .CLK(clk), .Q(arr[444]) );
  DFFPOSX1 arr_reg_13__14_ ( .D(n7201), .CLK(clk), .Q(arr[443]) );
  DFFPOSX1 arr_reg_13__13_ ( .D(n7200), .CLK(clk), .Q(arr[442]) );
  DFFPOSX1 arr_reg_13__12_ ( .D(n7199), .CLK(clk), .Q(arr[441]) );
  DFFPOSX1 arr_reg_13__11_ ( .D(n7198), .CLK(clk), .Q(arr[440]) );
  DFFPOSX1 arr_reg_13__10_ ( .D(n7197), .CLK(clk), .Q(arr[439]) );
  DFFPOSX1 arr_reg_13__9_ ( .D(n7196), .CLK(clk), .Q(arr[438]) );
  DFFPOSX1 arr_reg_13__8_ ( .D(n7195), .CLK(clk), .Q(arr[437]) );
  DFFPOSX1 arr_reg_13__7_ ( .D(n7194), .CLK(clk), .Q(arr[436]) );
  DFFPOSX1 arr_reg_13__6_ ( .D(n7193), .CLK(clk), .Q(arr[435]) );
  DFFPOSX1 arr_reg_13__5_ ( .D(n7192), .CLK(clk), .Q(arr[434]) );
  DFFPOSX1 arr_reg_13__4_ ( .D(n7191), .CLK(clk), .Q(arr[433]) );
  DFFPOSX1 arr_reg_13__3_ ( .D(n7190), .CLK(clk), .Q(arr[432]) );
  DFFPOSX1 arr_reg_13__2_ ( .D(n7189), .CLK(clk), .Q(arr[431]) );
  DFFPOSX1 arr_reg_13__1_ ( .D(n7188), .CLK(clk), .Q(arr[430]) );
  DFFPOSX1 arr_reg_13__0_ ( .D(n7187), .CLK(clk), .Q(arr[429]) );
  DFFPOSX1 arr_reg_12__32_ ( .D(n7186), .CLK(clk), .Q(arr[428]) );
  DFFPOSX1 arr_reg_12__31_ ( .D(n7185), .CLK(clk), .Q(arr[427]) );
  DFFPOSX1 arr_reg_12__30_ ( .D(n7184), .CLK(clk), .Q(arr[426]) );
  DFFPOSX1 arr_reg_12__29_ ( .D(n7183), .CLK(clk), .Q(arr[425]) );
  DFFPOSX1 arr_reg_12__28_ ( .D(n7182), .CLK(clk), .Q(arr[424]) );
  DFFPOSX1 arr_reg_12__27_ ( .D(n7181), .CLK(clk), .Q(arr[423]) );
  DFFPOSX1 arr_reg_12__26_ ( .D(n7180), .CLK(clk), .Q(arr[422]) );
  DFFPOSX1 arr_reg_12__25_ ( .D(n7179), .CLK(clk), .Q(arr[421]) );
  DFFPOSX1 arr_reg_12__24_ ( .D(n7178), .CLK(clk), .Q(arr[420]) );
  DFFPOSX1 arr_reg_12__23_ ( .D(n7177), .CLK(clk), .Q(arr[419]) );
  DFFPOSX1 arr_reg_12__22_ ( .D(n7176), .CLK(clk), .Q(arr[418]) );
  DFFPOSX1 arr_reg_12__21_ ( .D(n7175), .CLK(clk), .Q(arr[417]) );
  DFFPOSX1 arr_reg_12__20_ ( .D(n7174), .CLK(clk), .Q(arr[416]) );
  DFFPOSX1 arr_reg_12__19_ ( .D(n7173), .CLK(clk), .Q(arr[415]) );
  DFFPOSX1 arr_reg_12__18_ ( .D(n7172), .CLK(clk), .Q(arr[414]) );
  DFFPOSX1 arr_reg_12__17_ ( .D(n7171), .CLK(clk), .Q(arr[413]) );
  DFFPOSX1 arr_reg_12__16_ ( .D(n7170), .CLK(clk), .Q(arr[412]) );
  DFFPOSX1 arr_reg_12__15_ ( .D(n7169), .CLK(clk), .Q(arr[411]) );
  DFFPOSX1 arr_reg_12__14_ ( .D(n7168), .CLK(clk), .Q(arr[410]) );
  DFFPOSX1 arr_reg_12__13_ ( .D(n7167), .CLK(clk), .Q(arr[409]) );
  DFFPOSX1 arr_reg_12__12_ ( .D(n7166), .CLK(clk), .Q(arr[408]) );
  DFFPOSX1 arr_reg_12__11_ ( .D(n7165), .CLK(clk), .Q(arr[407]) );
  DFFPOSX1 arr_reg_12__10_ ( .D(n7164), .CLK(clk), .Q(arr[406]) );
  DFFPOSX1 arr_reg_12__9_ ( .D(n7163), .CLK(clk), .Q(arr[405]) );
  DFFPOSX1 arr_reg_12__8_ ( .D(n7162), .CLK(clk), .Q(arr[404]) );
  DFFPOSX1 arr_reg_12__7_ ( .D(n7161), .CLK(clk), .Q(arr[403]) );
  DFFPOSX1 arr_reg_12__6_ ( .D(n7160), .CLK(clk), .Q(arr[402]) );
  DFFPOSX1 arr_reg_12__5_ ( .D(n7159), .CLK(clk), .Q(arr[401]) );
  DFFPOSX1 arr_reg_12__4_ ( .D(n7158), .CLK(clk), .Q(arr[400]) );
  DFFPOSX1 arr_reg_12__3_ ( .D(n7157), .CLK(clk), .Q(arr[399]) );
  DFFPOSX1 arr_reg_12__2_ ( .D(n7156), .CLK(clk), .Q(arr[398]) );
  DFFPOSX1 arr_reg_12__1_ ( .D(n7155), .CLK(clk), .Q(arr[397]) );
  DFFPOSX1 arr_reg_12__0_ ( .D(n7154), .CLK(clk), .Q(arr[396]) );
  DFFPOSX1 arr_reg_11__32_ ( .D(n7153), .CLK(clk), .Q(arr[395]) );
  DFFPOSX1 arr_reg_11__31_ ( .D(n7152), .CLK(clk), .Q(arr[394]) );
  DFFPOSX1 arr_reg_11__30_ ( .D(n7151), .CLK(clk), .Q(arr[393]) );
  DFFPOSX1 arr_reg_11__29_ ( .D(n7150), .CLK(clk), .Q(arr[392]) );
  DFFPOSX1 arr_reg_11__28_ ( .D(n7149), .CLK(clk), .Q(arr[391]) );
  DFFPOSX1 arr_reg_11__27_ ( .D(n7148), .CLK(clk), .Q(arr[390]) );
  DFFPOSX1 arr_reg_11__26_ ( .D(n7147), .CLK(clk), .Q(arr[389]) );
  DFFPOSX1 arr_reg_11__25_ ( .D(n7146), .CLK(clk), .Q(arr[388]) );
  DFFPOSX1 arr_reg_11__24_ ( .D(n7145), .CLK(clk), .Q(arr[387]) );
  DFFPOSX1 arr_reg_11__23_ ( .D(n7144), .CLK(clk), .Q(arr[386]) );
  DFFPOSX1 arr_reg_11__22_ ( .D(n7143), .CLK(clk), .Q(arr[385]) );
  DFFPOSX1 arr_reg_11__21_ ( .D(n7142), .CLK(clk), .Q(arr[384]) );
  DFFPOSX1 arr_reg_11__20_ ( .D(n7141), .CLK(clk), .Q(arr[383]) );
  DFFPOSX1 arr_reg_11__19_ ( .D(n7140), .CLK(clk), .Q(arr[382]) );
  DFFPOSX1 arr_reg_11__18_ ( .D(n7139), .CLK(clk), .Q(arr[381]) );
  DFFPOSX1 arr_reg_11__17_ ( .D(n7138), .CLK(clk), .Q(arr[380]) );
  DFFPOSX1 arr_reg_11__16_ ( .D(n7137), .CLK(clk), .Q(arr[379]) );
  DFFPOSX1 arr_reg_11__15_ ( .D(n7136), .CLK(clk), .Q(arr[378]) );
  DFFPOSX1 arr_reg_11__14_ ( .D(n7135), .CLK(clk), .Q(arr[377]) );
  DFFPOSX1 arr_reg_11__13_ ( .D(n7134), .CLK(clk), .Q(arr[376]) );
  DFFPOSX1 arr_reg_11__12_ ( .D(n7133), .CLK(clk), .Q(arr[375]) );
  DFFPOSX1 arr_reg_11__11_ ( .D(n7132), .CLK(clk), .Q(arr[374]) );
  DFFPOSX1 arr_reg_11__10_ ( .D(n7131), .CLK(clk), .Q(arr[373]) );
  DFFPOSX1 arr_reg_11__9_ ( .D(n7130), .CLK(clk), .Q(arr[372]) );
  DFFPOSX1 arr_reg_11__8_ ( .D(n7129), .CLK(clk), .Q(arr[371]) );
  DFFPOSX1 arr_reg_11__7_ ( .D(n7128), .CLK(clk), .Q(arr[370]) );
  DFFPOSX1 arr_reg_11__6_ ( .D(n7127), .CLK(clk), .Q(arr[369]) );
  DFFPOSX1 arr_reg_11__5_ ( .D(n7126), .CLK(clk), .Q(arr[368]) );
  DFFPOSX1 arr_reg_11__4_ ( .D(n7125), .CLK(clk), .Q(arr[367]) );
  DFFPOSX1 arr_reg_11__3_ ( .D(n7124), .CLK(clk), .Q(arr[366]) );
  DFFPOSX1 arr_reg_11__2_ ( .D(n7123), .CLK(clk), .Q(arr[365]) );
  DFFPOSX1 arr_reg_11__1_ ( .D(n7122), .CLK(clk), .Q(arr[364]) );
  DFFPOSX1 arr_reg_11__0_ ( .D(n7121), .CLK(clk), .Q(arr[363]) );
  DFFPOSX1 arr_reg_10__32_ ( .D(n7120), .CLK(clk), .Q(arr[362]) );
  DFFPOSX1 arr_reg_10__31_ ( .D(n7119), .CLK(clk), .Q(arr[361]) );
  DFFPOSX1 arr_reg_10__30_ ( .D(n7118), .CLK(clk), .Q(arr[360]) );
  DFFPOSX1 arr_reg_10__29_ ( .D(n7117), .CLK(clk), .Q(arr[359]) );
  DFFPOSX1 arr_reg_10__28_ ( .D(n7116), .CLK(clk), .Q(arr[358]) );
  DFFPOSX1 arr_reg_10__27_ ( .D(n7115), .CLK(clk), .Q(arr[357]) );
  DFFPOSX1 arr_reg_10__26_ ( .D(n7114), .CLK(clk), .Q(arr[356]) );
  DFFPOSX1 arr_reg_10__25_ ( .D(n7113), .CLK(clk), .Q(arr[355]) );
  DFFPOSX1 arr_reg_10__24_ ( .D(n7112), .CLK(clk), .Q(arr[354]) );
  DFFPOSX1 arr_reg_10__23_ ( .D(n7111), .CLK(clk), .Q(arr[353]) );
  DFFPOSX1 arr_reg_10__22_ ( .D(n7110), .CLK(clk), .Q(arr[352]) );
  DFFPOSX1 arr_reg_10__21_ ( .D(n7109), .CLK(clk), .Q(arr[351]) );
  DFFPOSX1 arr_reg_10__20_ ( .D(n7108), .CLK(clk), .Q(arr[350]) );
  DFFPOSX1 arr_reg_10__19_ ( .D(n7107), .CLK(clk), .Q(arr[349]) );
  DFFPOSX1 arr_reg_10__18_ ( .D(n7106), .CLK(clk), .Q(arr[348]) );
  DFFPOSX1 arr_reg_10__17_ ( .D(n7105), .CLK(clk), .Q(arr[347]) );
  DFFPOSX1 arr_reg_10__16_ ( .D(n7104), .CLK(clk), .Q(arr[346]) );
  DFFPOSX1 arr_reg_10__15_ ( .D(n7103), .CLK(clk), .Q(arr[345]) );
  DFFPOSX1 arr_reg_10__14_ ( .D(n7102), .CLK(clk), .Q(arr[344]) );
  DFFPOSX1 arr_reg_10__13_ ( .D(n7101), .CLK(clk), .Q(arr[343]) );
  DFFPOSX1 arr_reg_10__12_ ( .D(n7100), .CLK(clk), .Q(arr[342]) );
  DFFPOSX1 arr_reg_10__11_ ( .D(n7099), .CLK(clk), .Q(arr[341]) );
  DFFPOSX1 arr_reg_10__10_ ( .D(n7098), .CLK(clk), .Q(arr[340]) );
  DFFPOSX1 arr_reg_10__9_ ( .D(n7097), .CLK(clk), .Q(arr[339]) );
  DFFPOSX1 arr_reg_10__8_ ( .D(n7096), .CLK(clk), .Q(arr[338]) );
  DFFPOSX1 arr_reg_10__7_ ( .D(n7095), .CLK(clk), .Q(arr[337]) );
  DFFPOSX1 arr_reg_10__6_ ( .D(n7094), .CLK(clk), .Q(arr[336]) );
  DFFPOSX1 arr_reg_10__5_ ( .D(n7093), .CLK(clk), .Q(arr[335]) );
  DFFPOSX1 arr_reg_10__4_ ( .D(n7092), .CLK(clk), .Q(arr[334]) );
  DFFPOSX1 arr_reg_10__3_ ( .D(n7091), .CLK(clk), .Q(arr[333]) );
  DFFPOSX1 arr_reg_10__2_ ( .D(n7090), .CLK(clk), .Q(arr[332]) );
  DFFPOSX1 arr_reg_10__1_ ( .D(n7089), .CLK(clk), .Q(arr[331]) );
  DFFPOSX1 arr_reg_10__0_ ( .D(n7088), .CLK(clk), .Q(arr[330]) );
  DFFPOSX1 arr_reg_9__32_ ( .D(n7087), .CLK(clk), .Q(arr[329]) );
  DFFPOSX1 arr_reg_9__31_ ( .D(n7086), .CLK(clk), .Q(arr[328]) );
  DFFPOSX1 arr_reg_9__30_ ( .D(n7085), .CLK(clk), .Q(arr[327]) );
  DFFPOSX1 arr_reg_9__29_ ( .D(n7084), .CLK(clk), .Q(arr[326]) );
  DFFPOSX1 arr_reg_9__28_ ( .D(n7083), .CLK(clk), .Q(arr[325]) );
  DFFPOSX1 arr_reg_9__27_ ( .D(n7082), .CLK(clk), .Q(arr[324]) );
  DFFPOSX1 arr_reg_9__26_ ( .D(n7081), .CLK(clk), .Q(arr[323]) );
  DFFPOSX1 arr_reg_9__25_ ( .D(n7080), .CLK(clk), .Q(arr[322]) );
  DFFPOSX1 arr_reg_9__24_ ( .D(n7079), .CLK(clk), .Q(arr[321]) );
  DFFPOSX1 arr_reg_9__23_ ( .D(n7078), .CLK(clk), .Q(arr[320]) );
  DFFPOSX1 arr_reg_9__22_ ( .D(n7077), .CLK(clk), .Q(arr[319]) );
  DFFPOSX1 arr_reg_9__21_ ( .D(n7076), .CLK(clk), .Q(arr[318]) );
  DFFPOSX1 arr_reg_9__20_ ( .D(n7075), .CLK(clk), .Q(arr[317]) );
  DFFPOSX1 arr_reg_9__19_ ( .D(n7074), .CLK(clk), .Q(arr[316]) );
  DFFPOSX1 arr_reg_9__18_ ( .D(n7073), .CLK(clk), .Q(arr[315]) );
  DFFPOSX1 arr_reg_9__17_ ( .D(n7072), .CLK(clk), .Q(arr[314]) );
  DFFPOSX1 arr_reg_9__16_ ( .D(n7071), .CLK(clk), .Q(arr[313]) );
  DFFPOSX1 arr_reg_9__15_ ( .D(n7070), .CLK(clk), .Q(arr[312]) );
  DFFPOSX1 arr_reg_9__14_ ( .D(n7069), .CLK(clk), .Q(arr[311]) );
  DFFPOSX1 arr_reg_9__13_ ( .D(n7068), .CLK(clk), .Q(arr[310]) );
  DFFPOSX1 arr_reg_9__12_ ( .D(n7067), .CLK(clk), .Q(arr[309]) );
  DFFPOSX1 arr_reg_9__11_ ( .D(n7066), .CLK(clk), .Q(arr[308]) );
  DFFPOSX1 arr_reg_9__10_ ( .D(n7065), .CLK(clk), .Q(arr[307]) );
  DFFPOSX1 arr_reg_9__9_ ( .D(n7064), .CLK(clk), .Q(arr[306]) );
  DFFPOSX1 arr_reg_9__8_ ( .D(n7063), .CLK(clk), .Q(arr[305]) );
  DFFPOSX1 arr_reg_9__7_ ( .D(n7062), .CLK(clk), .Q(arr[304]) );
  DFFPOSX1 arr_reg_9__6_ ( .D(n7061), .CLK(clk), .Q(arr[303]) );
  DFFPOSX1 arr_reg_9__5_ ( .D(n7060), .CLK(clk), .Q(arr[302]) );
  DFFPOSX1 arr_reg_9__4_ ( .D(n7059), .CLK(clk), .Q(arr[301]) );
  DFFPOSX1 arr_reg_9__3_ ( .D(n7058), .CLK(clk), .Q(arr[300]) );
  DFFPOSX1 arr_reg_9__2_ ( .D(n7057), .CLK(clk), .Q(arr[299]) );
  DFFPOSX1 arr_reg_9__1_ ( .D(n7056), .CLK(clk), .Q(arr[298]) );
  DFFPOSX1 arr_reg_9__0_ ( .D(n7055), .CLK(clk), .Q(arr[297]) );
  DFFPOSX1 arr_reg_8__32_ ( .D(n7054), .CLK(clk), .Q(arr[296]) );
  DFFPOSX1 arr_reg_8__31_ ( .D(n7053), .CLK(clk), .Q(arr[295]) );
  DFFPOSX1 arr_reg_8__30_ ( .D(n7052), .CLK(clk), .Q(arr[294]) );
  DFFPOSX1 arr_reg_8__29_ ( .D(n7051), .CLK(clk), .Q(arr[293]) );
  DFFPOSX1 arr_reg_8__28_ ( .D(n7050), .CLK(clk), .Q(arr[292]) );
  DFFPOSX1 arr_reg_8__27_ ( .D(n7049), .CLK(clk), .Q(arr[291]) );
  DFFPOSX1 arr_reg_8__26_ ( .D(n7048), .CLK(clk), .Q(arr[290]) );
  DFFPOSX1 arr_reg_8__25_ ( .D(n7047), .CLK(clk), .Q(arr[289]) );
  DFFPOSX1 arr_reg_8__24_ ( .D(n7046), .CLK(clk), .Q(arr[288]) );
  DFFPOSX1 arr_reg_8__23_ ( .D(n7045), .CLK(clk), .Q(arr[287]) );
  DFFPOSX1 arr_reg_8__22_ ( .D(n7044), .CLK(clk), .Q(arr[286]) );
  DFFPOSX1 arr_reg_8__21_ ( .D(n7043), .CLK(clk), .Q(arr[285]) );
  DFFPOSX1 arr_reg_8__20_ ( .D(n7042), .CLK(clk), .Q(arr[284]) );
  DFFPOSX1 arr_reg_8__19_ ( .D(n7041), .CLK(clk), .Q(arr[283]) );
  DFFPOSX1 arr_reg_8__18_ ( .D(n7040), .CLK(clk), .Q(arr[282]) );
  DFFPOSX1 arr_reg_8__17_ ( .D(n7039), .CLK(clk), .Q(arr[281]) );
  DFFPOSX1 arr_reg_8__16_ ( .D(n7038), .CLK(clk), .Q(arr[280]) );
  DFFPOSX1 arr_reg_8__15_ ( .D(n7037), .CLK(clk), .Q(arr[279]) );
  DFFPOSX1 arr_reg_8__14_ ( .D(n7036), .CLK(clk), .Q(arr[278]) );
  DFFPOSX1 arr_reg_8__13_ ( .D(n7035), .CLK(clk), .Q(arr[277]) );
  DFFPOSX1 arr_reg_8__12_ ( .D(n7034), .CLK(clk), .Q(arr[276]) );
  DFFPOSX1 arr_reg_8__11_ ( .D(n7033), .CLK(clk), .Q(arr[275]) );
  DFFPOSX1 arr_reg_8__10_ ( .D(n7032), .CLK(clk), .Q(arr[274]) );
  DFFPOSX1 arr_reg_8__9_ ( .D(n7031), .CLK(clk), .Q(arr[273]) );
  DFFPOSX1 arr_reg_8__8_ ( .D(n7030), .CLK(clk), .Q(arr[272]) );
  DFFPOSX1 arr_reg_8__7_ ( .D(n7029), .CLK(clk), .Q(arr[271]) );
  DFFPOSX1 arr_reg_8__6_ ( .D(n7028), .CLK(clk), .Q(arr[270]) );
  DFFPOSX1 arr_reg_8__5_ ( .D(n7027), .CLK(clk), .Q(arr[269]) );
  DFFPOSX1 arr_reg_8__4_ ( .D(n7026), .CLK(clk), .Q(arr[268]) );
  DFFPOSX1 arr_reg_8__3_ ( .D(n7025), .CLK(clk), .Q(arr[267]) );
  DFFPOSX1 arr_reg_8__2_ ( .D(n7024), .CLK(clk), .Q(arr[266]) );
  DFFPOSX1 arr_reg_8__1_ ( .D(n7023), .CLK(clk), .Q(arr[265]) );
  DFFPOSX1 arr_reg_8__0_ ( .D(n7022), .CLK(clk), .Q(arr[264]) );
  DFFPOSX1 arr_reg_7__32_ ( .D(n7021), .CLK(clk), .Q(arr[263]) );
  DFFPOSX1 arr_reg_7__31_ ( .D(n7020), .CLK(clk), .Q(arr[262]) );
  DFFPOSX1 arr_reg_7__30_ ( .D(n7019), .CLK(clk), .Q(arr[261]) );
  DFFPOSX1 arr_reg_7__29_ ( .D(n7018), .CLK(clk), .Q(arr[260]) );
  DFFPOSX1 arr_reg_7__28_ ( .D(n7017), .CLK(clk), .Q(arr[259]) );
  DFFPOSX1 arr_reg_7__27_ ( .D(n7016), .CLK(clk), .Q(arr[258]) );
  DFFPOSX1 arr_reg_7__26_ ( .D(n7015), .CLK(clk), .Q(arr[257]) );
  DFFPOSX1 arr_reg_7__25_ ( .D(n7014), .CLK(clk), .Q(arr[256]) );
  DFFPOSX1 arr_reg_7__24_ ( .D(n7013), .CLK(clk), .Q(arr[255]) );
  DFFPOSX1 arr_reg_7__23_ ( .D(n7012), .CLK(clk), .Q(arr[254]) );
  DFFPOSX1 arr_reg_7__22_ ( .D(n7011), .CLK(clk), .Q(arr[253]) );
  DFFPOSX1 arr_reg_7__21_ ( .D(n7010), .CLK(clk), .Q(arr[252]) );
  DFFPOSX1 arr_reg_7__20_ ( .D(n7009), .CLK(clk), .Q(arr[251]) );
  DFFPOSX1 arr_reg_7__19_ ( .D(n7008), .CLK(clk), .Q(arr[250]) );
  DFFPOSX1 arr_reg_7__18_ ( .D(n7007), .CLK(clk), .Q(arr[249]) );
  DFFPOSX1 arr_reg_7__17_ ( .D(n7006), .CLK(clk), .Q(arr[248]) );
  DFFPOSX1 arr_reg_7__16_ ( .D(n7005), .CLK(clk), .Q(arr[247]) );
  DFFPOSX1 arr_reg_7__15_ ( .D(n7004), .CLK(clk), .Q(arr[246]) );
  DFFPOSX1 arr_reg_7__14_ ( .D(n7003), .CLK(clk), .Q(arr[245]) );
  DFFPOSX1 arr_reg_7__13_ ( .D(n7002), .CLK(clk), .Q(arr[244]) );
  DFFPOSX1 arr_reg_7__12_ ( .D(n7001), .CLK(clk), .Q(arr[243]) );
  DFFPOSX1 arr_reg_7__11_ ( .D(n7000), .CLK(clk), .Q(arr[242]) );
  DFFPOSX1 arr_reg_7__10_ ( .D(n6999), .CLK(clk), .Q(arr[241]) );
  DFFPOSX1 arr_reg_7__9_ ( .D(n6998), .CLK(clk), .Q(arr[240]) );
  DFFPOSX1 arr_reg_7__8_ ( .D(n6997), .CLK(clk), .Q(arr[239]) );
  DFFPOSX1 arr_reg_7__7_ ( .D(n6996), .CLK(clk), .Q(arr[238]) );
  DFFPOSX1 arr_reg_7__6_ ( .D(n6995), .CLK(clk), .Q(arr[237]) );
  DFFPOSX1 arr_reg_7__5_ ( .D(n6994), .CLK(clk), .Q(arr[236]) );
  DFFPOSX1 arr_reg_7__4_ ( .D(n6993), .CLK(clk), .Q(arr[235]) );
  DFFPOSX1 arr_reg_7__3_ ( .D(n6992), .CLK(clk), .Q(arr[234]) );
  DFFPOSX1 arr_reg_7__2_ ( .D(n6991), .CLK(clk), .Q(arr[233]) );
  DFFPOSX1 arr_reg_7__1_ ( .D(n6990), .CLK(clk), .Q(arr[232]) );
  DFFPOSX1 arr_reg_7__0_ ( .D(n6989), .CLK(clk), .Q(arr[231]) );
  DFFPOSX1 arr_reg_6__32_ ( .D(n6988), .CLK(clk), .Q(arr[230]) );
  DFFPOSX1 arr_reg_6__31_ ( .D(n6987), .CLK(clk), .Q(arr[229]) );
  DFFPOSX1 arr_reg_6__30_ ( .D(n6986), .CLK(clk), .Q(arr[228]) );
  DFFPOSX1 arr_reg_6__29_ ( .D(n6985), .CLK(clk), .Q(arr[227]) );
  DFFPOSX1 arr_reg_6__28_ ( .D(n6984), .CLK(clk), .Q(arr[226]) );
  DFFPOSX1 arr_reg_6__27_ ( .D(n6983), .CLK(clk), .Q(arr[225]) );
  DFFPOSX1 arr_reg_6__26_ ( .D(n6982), .CLK(clk), .Q(arr[224]) );
  DFFPOSX1 arr_reg_6__25_ ( .D(n6981), .CLK(clk), .Q(arr[223]) );
  DFFPOSX1 arr_reg_6__24_ ( .D(n6980), .CLK(clk), .Q(arr[222]) );
  DFFPOSX1 arr_reg_6__23_ ( .D(n6979), .CLK(clk), .Q(arr[221]) );
  DFFPOSX1 arr_reg_6__22_ ( .D(n6978), .CLK(clk), .Q(arr[220]) );
  DFFPOSX1 arr_reg_6__21_ ( .D(n6977), .CLK(clk), .Q(arr[219]) );
  DFFPOSX1 arr_reg_6__20_ ( .D(n6976), .CLK(clk), .Q(arr[218]) );
  DFFPOSX1 arr_reg_6__19_ ( .D(n6975), .CLK(clk), .Q(arr[217]) );
  DFFPOSX1 arr_reg_6__18_ ( .D(n6974), .CLK(clk), .Q(arr[216]) );
  DFFPOSX1 arr_reg_6__17_ ( .D(n6973), .CLK(clk), .Q(arr[215]) );
  DFFPOSX1 arr_reg_6__16_ ( .D(n6972), .CLK(clk), .Q(arr[214]) );
  DFFPOSX1 arr_reg_6__15_ ( .D(n6971), .CLK(clk), .Q(arr[213]) );
  DFFPOSX1 arr_reg_6__14_ ( .D(n6970), .CLK(clk), .Q(arr[212]) );
  DFFPOSX1 arr_reg_6__13_ ( .D(n6969), .CLK(clk), .Q(arr[211]) );
  DFFPOSX1 arr_reg_6__12_ ( .D(n6968), .CLK(clk), .Q(arr[210]) );
  DFFPOSX1 arr_reg_6__11_ ( .D(n6967), .CLK(clk), .Q(arr[209]) );
  DFFPOSX1 arr_reg_6__10_ ( .D(n6966), .CLK(clk), .Q(arr[208]) );
  DFFPOSX1 arr_reg_6__9_ ( .D(n6965), .CLK(clk), .Q(arr[207]) );
  DFFPOSX1 arr_reg_6__8_ ( .D(n6964), .CLK(clk), .Q(arr[206]) );
  DFFPOSX1 arr_reg_6__7_ ( .D(n6963), .CLK(clk), .Q(arr[205]) );
  DFFPOSX1 arr_reg_6__6_ ( .D(n6962), .CLK(clk), .Q(arr[204]) );
  DFFPOSX1 arr_reg_6__5_ ( .D(n6961), .CLK(clk), .Q(arr[203]) );
  DFFPOSX1 arr_reg_6__4_ ( .D(n6960), .CLK(clk), .Q(arr[202]) );
  DFFPOSX1 arr_reg_6__3_ ( .D(n6959), .CLK(clk), .Q(arr[201]) );
  DFFPOSX1 arr_reg_6__2_ ( .D(n6958), .CLK(clk), .Q(arr[200]) );
  DFFPOSX1 arr_reg_6__1_ ( .D(n6957), .CLK(clk), .Q(arr[199]) );
  DFFPOSX1 arr_reg_6__0_ ( .D(n6956), .CLK(clk), .Q(arr[198]) );
  DFFPOSX1 arr_reg_5__32_ ( .D(n6955), .CLK(clk), .Q(arr[197]) );
  DFFPOSX1 arr_reg_5__31_ ( .D(n6954), .CLK(clk), .Q(arr[196]) );
  DFFPOSX1 arr_reg_5__30_ ( .D(n6953), .CLK(clk), .Q(arr[195]) );
  DFFPOSX1 arr_reg_5__29_ ( .D(n6952), .CLK(clk), .Q(arr[194]) );
  DFFPOSX1 arr_reg_5__28_ ( .D(n6951), .CLK(clk), .Q(arr[193]) );
  DFFPOSX1 arr_reg_5__27_ ( .D(n6950), .CLK(clk), .Q(arr[192]) );
  DFFPOSX1 arr_reg_5__26_ ( .D(n6949), .CLK(clk), .Q(arr[191]) );
  DFFPOSX1 arr_reg_5__25_ ( .D(n6948), .CLK(clk), .Q(arr[190]) );
  DFFPOSX1 arr_reg_5__24_ ( .D(n6947), .CLK(clk), .Q(arr[189]) );
  DFFPOSX1 arr_reg_5__23_ ( .D(n6946), .CLK(clk), .Q(arr[188]) );
  DFFPOSX1 arr_reg_5__22_ ( .D(n6945), .CLK(clk), .Q(arr[187]) );
  DFFPOSX1 arr_reg_5__21_ ( .D(n6944), .CLK(clk), .Q(arr[186]) );
  DFFPOSX1 arr_reg_5__20_ ( .D(n6943), .CLK(clk), .Q(arr[185]) );
  DFFPOSX1 arr_reg_5__19_ ( .D(n6942), .CLK(clk), .Q(arr[184]) );
  DFFPOSX1 arr_reg_5__18_ ( .D(n6941), .CLK(clk), .Q(arr[183]) );
  DFFPOSX1 arr_reg_5__17_ ( .D(n6940), .CLK(clk), .Q(arr[182]) );
  DFFPOSX1 arr_reg_5__16_ ( .D(n6939), .CLK(clk), .Q(arr[181]) );
  DFFPOSX1 arr_reg_5__15_ ( .D(n6938), .CLK(clk), .Q(arr[180]) );
  DFFPOSX1 arr_reg_5__14_ ( .D(n6937), .CLK(clk), .Q(arr[179]) );
  DFFPOSX1 arr_reg_5__13_ ( .D(n6936), .CLK(clk), .Q(arr[178]) );
  DFFPOSX1 arr_reg_5__12_ ( .D(n6935), .CLK(clk), .Q(arr[177]) );
  DFFPOSX1 arr_reg_5__11_ ( .D(n6934), .CLK(clk), .Q(arr[176]) );
  DFFPOSX1 arr_reg_5__10_ ( .D(n6933), .CLK(clk), .Q(arr[175]) );
  DFFPOSX1 arr_reg_5__9_ ( .D(n6932), .CLK(clk), .Q(arr[174]) );
  DFFPOSX1 arr_reg_5__8_ ( .D(n6931), .CLK(clk), .Q(arr[173]) );
  DFFPOSX1 arr_reg_5__7_ ( .D(n6930), .CLK(clk), .Q(arr[172]) );
  DFFPOSX1 arr_reg_5__6_ ( .D(n6929), .CLK(clk), .Q(arr[171]) );
  DFFPOSX1 arr_reg_5__5_ ( .D(n6928), .CLK(clk), .Q(arr[170]) );
  DFFPOSX1 arr_reg_5__4_ ( .D(n6927), .CLK(clk), .Q(arr[169]) );
  DFFPOSX1 arr_reg_5__3_ ( .D(n6926), .CLK(clk), .Q(arr[168]) );
  DFFPOSX1 arr_reg_5__2_ ( .D(n6925), .CLK(clk), .Q(arr[167]) );
  DFFPOSX1 arr_reg_5__1_ ( .D(n6924), .CLK(clk), .Q(arr[166]) );
  DFFPOSX1 arr_reg_5__0_ ( .D(n6923), .CLK(clk), .Q(arr[165]) );
  DFFPOSX1 arr_reg_4__32_ ( .D(n6922), .CLK(clk), .Q(arr[164]) );
  DFFPOSX1 arr_reg_4__31_ ( .D(n6921), .CLK(clk), .Q(arr[163]) );
  DFFPOSX1 arr_reg_4__30_ ( .D(n6920), .CLK(clk), .Q(arr[162]) );
  DFFPOSX1 arr_reg_4__29_ ( .D(n6919), .CLK(clk), .Q(arr[161]) );
  DFFPOSX1 arr_reg_4__28_ ( .D(n6918), .CLK(clk), .Q(arr[160]) );
  DFFPOSX1 arr_reg_4__27_ ( .D(n6917), .CLK(clk), .Q(arr[159]) );
  DFFPOSX1 arr_reg_4__26_ ( .D(n6916), .CLK(clk), .Q(arr[158]) );
  DFFPOSX1 arr_reg_4__25_ ( .D(n6915), .CLK(clk), .Q(arr[157]) );
  DFFPOSX1 arr_reg_4__24_ ( .D(n6914), .CLK(clk), .Q(arr[156]) );
  DFFPOSX1 arr_reg_4__23_ ( .D(n6913), .CLK(clk), .Q(arr[155]) );
  DFFPOSX1 arr_reg_4__22_ ( .D(n6912), .CLK(clk), .Q(arr[154]) );
  DFFPOSX1 arr_reg_4__21_ ( .D(n6911), .CLK(clk), .Q(arr[153]) );
  DFFPOSX1 arr_reg_4__20_ ( .D(n6910), .CLK(clk), .Q(arr[152]) );
  DFFPOSX1 arr_reg_4__19_ ( .D(n6909), .CLK(clk), .Q(arr[151]) );
  DFFPOSX1 arr_reg_4__18_ ( .D(n6908), .CLK(clk), .Q(arr[150]) );
  DFFPOSX1 arr_reg_4__17_ ( .D(n6907), .CLK(clk), .Q(arr[149]) );
  DFFPOSX1 arr_reg_4__16_ ( .D(n6906), .CLK(clk), .Q(arr[148]) );
  DFFPOSX1 arr_reg_4__15_ ( .D(n6905), .CLK(clk), .Q(arr[147]) );
  DFFPOSX1 arr_reg_4__14_ ( .D(n6904), .CLK(clk), .Q(arr[146]) );
  DFFPOSX1 arr_reg_4__13_ ( .D(n6903), .CLK(clk), .Q(arr[145]) );
  DFFPOSX1 arr_reg_4__12_ ( .D(n6902), .CLK(clk), .Q(arr[144]) );
  DFFPOSX1 arr_reg_4__11_ ( .D(n6901), .CLK(clk), .Q(arr[143]) );
  DFFPOSX1 arr_reg_4__10_ ( .D(n6900), .CLK(clk), .Q(arr[142]) );
  DFFPOSX1 arr_reg_4__9_ ( .D(n6899), .CLK(clk), .Q(arr[141]) );
  DFFPOSX1 arr_reg_4__8_ ( .D(n6898), .CLK(clk), .Q(arr[140]) );
  DFFPOSX1 arr_reg_4__7_ ( .D(n6897), .CLK(clk), .Q(arr[139]) );
  DFFPOSX1 arr_reg_4__6_ ( .D(n6896), .CLK(clk), .Q(arr[138]) );
  DFFPOSX1 arr_reg_4__5_ ( .D(n6895), .CLK(clk), .Q(arr[137]) );
  DFFPOSX1 arr_reg_4__4_ ( .D(n6894), .CLK(clk), .Q(arr[136]) );
  DFFPOSX1 arr_reg_4__3_ ( .D(n6893), .CLK(clk), .Q(arr[135]) );
  DFFPOSX1 arr_reg_4__2_ ( .D(n6892), .CLK(clk), .Q(arr[134]) );
  DFFPOSX1 arr_reg_4__1_ ( .D(n6891), .CLK(clk), .Q(arr[133]) );
  DFFPOSX1 arr_reg_4__0_ ( .D(n6890), .CLK(clk), .Q(arr[132]) );
  DFFPOSX1 arr_reg_3__32_ ( .D(n6889), .CLK(clk), .Q(arr[131]) );
  DFFPOSX1 arr_reg_3__31_ ( .D(n6888), .CLK(clk), .Q(arr[130]) );
  DFFPOSX1 arr_reg_3__30_ ( .D(n6887), .CLK(clk), .Q(arr[129]) );
  DFFPOSX1 arr_reg_3__29_ ( .D(n6886), .CLK(clk), .Q(arr[128]) );
  DFFPOSX1 arr_reg_3__28_ ( .D(n6885), .CLK(clk), .Q(arr[127]) );
  DFFPOSX1 arr_reg_3__27_ ( .D(n6884), .CLK(clk), .Q(arr[126]) );
  DFFPOSX1 arr_reg_3__26_ ( .D(n6883), .CLK(clk), .Q(arr[125]) );
  DFFPOSX1 arr_reg_3__25_ ( .D(n6882), .CLK(clk), .Q(arr[124]) );
  DFFPOSX1 arr_reg_3__24_ ( .D(n6881), .CLK(clk), .Q(arr[123]) );
  DFFPOSX1 arr_reg_3__23_ ( .D(n6880), .CLK(clk), .Q(arr[122]) );
  DFFPOSX1 arr_reg_3__22_ ( .D(n6879), .CLK(clk), .Q(arr[121]) );
  DFFPOSX1 arr_reg_3__21_ ( .D(n6878), .CLK(clk), .Q(arr[120]) );
  DFFPOSX1 arr_reg_3__20_ ( .D(n6877), .CLK(clk), .Q(arr[119]) );
  DFFPOSX1 arr_reg_3__19_ ( .D(n6876), .CLK(clk), .Q(arr[118]) );
  DFFPOSX1 arr_reg_3__18_ ( .D(n6875), .CLK(clk), .Q(arr[117]) );
  DFFPOSX1 arr_reg_3__17_ ( .D(n6874), .CLK(clk), .Q(arr[116]) );
  DFFPOSX1 arr_reg_3__16_ ( .D(n6873), .CLK(clk), .Q(arr[115]) );
  DFFPOSX1 arr_reg_3__15_ ( .D(n6872), .CLK(clk), .Q(arr[114]) );
  DFFPOSX1 arr_reg_3__14_ ( .D(n6871), .CLK(clk), .Q(arr[113]) );
  DFFPOSX1 arr_reg_3__13_ ( .D(n6870), .CLK(clk), .Q(arr[112]) );
  DFFPOSX1 arr_reg_3__12_ ( .D(n6869), .CLK(clk), .Q(arr[111]) );
  DFFPOSX1 arr_reg_3__11_ ( .D(n6868), .CLK(clk), .Q(arr[110]) );
  DFFPOSX1 arr_reg_3__10_ ( .D(n6867), .CLK(clk), .Q(arr[109]) );
  DFFPOSX1 arr_reg_3__9_ ( .D(n6866), .CLK(clk), .Q(arr[108]) );
  DFFPOSX1 arr_reg_3__8_ ( .D(n6865), .CLK(clk), .Q(arr[107]) );
  DFFPOSX1 arr_reg_3__7_ ( .D(n6864), .CLK(clk), .Q(arr[106]) );
  DFFPOSX1 arr_reg_3__6_ ( .D(n6863), .CLK(clk), .Q(arr[105]) );
  DFFPOSX1 arr_reg_3__5_ ( .D(n6862), .CLK(clk), .Q(arr[104]) );
  DFFPOSX1 arr_reg_3__4_ ( .D(n6861), .CLK(clk), .Q(arr[103]) );
  DFFPOSX1 arr_reg_3__3_ ( .D(n6860), .CLK(clk), .Q(arr[102]) );
  DFFPOSX1 arr_reg_3__2_ ( .D(n6859), .CLK(clk), .Q(arr[101]) );
  DFFPOSX1 arr_reg_3__1_ ( .D(n6858), .CLK(clk), .Q(arr[100]) );
  DFFPOSX1 arr_reg_3__0_ ( .D(n6857), .CLK(clk), .Q(arr[99]) );
  DFFPOSX1 arr_reg_2__32_ ( .D(n6856), .CLK(clk), .Q(arr[98]) );
  DFFPOSX1 arr_reg_2__31_ ( .D(n6855), .CLK(clk), .Q(arr[97]) );
  DFFPOSX1 arr_reg_2__30_ ( .D(n6854), .CLK(clk), .Q(arr[96]) );
  DFFPOSX1 arr_reg_2__29_ ( .D(n6853), .CLK(clk), .Q(arr[95]) );
  DFFPOSX1 arr_reg_2__28_ ( .D(n6852), .CLK(clk), .Q(arr[94]) );
  DFFPOSX1 arr_reg_2__27_ ( .D(n6851), .CLK(clk), .Q(arr[93]) );
  DFFPOSX1 arr_reg_2__26_ ( .D(n6850), .CLK(clk), .Q(arr[92]) );
  DFFPOSX1 arr_reg_2__25_ ( .D(n6849), .CLK(clk), .Q(arr[91]) );
  DFFPOSX1 arr_reg_2__24_ ( .D(n6848), .CLK(clk), .Q(arr[90]) );
  DFFPOSX1 arr_reg_2__23_ ( .D(n6847), .CLK(clk), .Q(arr[89]) );
  DFFPOSX1 arr_reg_2__22_ ( .D(n6846), .CLK(clk), .Q(arr[88]) );
  DFFPOSX1 arr_reg_2__21_ ( .D(n6845), .CLK(clk), .Q(arr[87]) );
  DFFPOSX1 arr_reg_2__20_ ( .D(n6844), .CLK(clk), .Q(arr[86]) );
  DFFPOSX1 arr_reg_2__19_ ( .D(n6843), .CLK(clk), .Q(arr[85]) );
  DFFPOSX1 arr_reg_2__18_ ( .D(n6842), .CLK(clk), .Q(arr[84]) );
  DFFPOSX1 arr_reg_2__17_ ( .D(n6841), .CLK(clk), .Q(arr[83]) );
  DFFPOSX1 arr_reg_2__16_ ( .D(n6840), .CLK(clk), .Q(arr[82]) );
  DFFPOSX1 arr_reg_2__15_ ( .D(n6839), .CLK(clk), .Q(arr[81]) );
  DFFPOSX1 arr_reg_2__14_ ( .D(n6838), .CLK(clk), .Q(arr[80]) );
  DFFPOSX1 arr_reg_2__13_ ( .D(n6837), .CLK(clk), .Q(arr[79]) );
  DFFPOSX1 arr_reg_2__12_ ( .D(n6836), .CLK(clk), .Q(arr[78]) );
  DFFPOSX1 arr_reg_2__11_ ( .D(n6835), .CLK(clk), .Q(arr[77]) );
  DFFPOSX1 arr_reg_2__10_ ( .D(n6834), .CLK(clk), .Q(arr[76]) );
  DFFPOSX1 arr_reg_2__9_ ( .D(n6833), .CLK(clk), .Q(arr[75]) );
  DFFPOSX1 arr_reg_2__8_ ( .D(n6832), .CLK(clk), .Q(arr[74]) );
  DFFPOSX1 arr_reg_2__7_ ( .D(n6831), .CLK(clk), .Q(arr[73]) );
  DFFPOSX1 arr_reg_2__6_ ( .D(n6830), .CLK(clk), .Q(arr[72]) );
  DFFPOSX1 arr_reg_2__5_ ( .D(n6829), .CLK(clk), .Q(arr[71]) );
  DFFPOSX1 arr_reg_2__4_ ( .D(n6828), .CLK(clk), .Q(arr[70]) );
  DFFPOSX1 arr_reg_2__3_ ( .D(n6827), .CLK(clk), .Q(arr[69]) );
  DFFPOSX1 arr_reg_2__2_ ( .D(n6826), .CLK(clk), .Q(arr[68]) );
  DFFPOSX1 arr_reg_2__1_ ( .D(n6825), .CLK(clk), .Q(arr[67]) );
  DFFPOSX1 arr_reg_2__0_ ( .D(n6824), .CLK(clk), .Q(arr[66]) );
  DFFPOSX1 arr_reg_1__32_ ( .D(n6823), .CLK(clk), .Q(arr[65]) );
  DFFPOSX1 arr_reg_1__31_ ( .D(n6822), .CLK(clk), .Q(arr[64]) );
  DFFPOSX1 arr_reg_1__30_ ( .D(n6821), .CLK(clk), .Q(arr[63]) );
  DFFPOSX1 arr_reg_1__29_ ( .D(n6820), .CLK(clk), .Q(arr[62]) );
  DFFPOSX1 arr_reg_1__28_ ( .D(n6819), .CLK(clk), .Q(arr[61]) );
  DFFPOSX1 arr_reg_1__27_ ( .D(n6818), .CLK(clk), .Q(arr[60]) );
  DFFPOSX1 arr_reg_1__26_ ( .D(n6817), .CLK(clk), .Q(arr[59]) );
  DFFPOSX1 arr_reg_1__25_ ( .D(n6816), .CLK(clk), .Q(arr[58]) );
  DFFPOSX1 arr_reg_1__24_ ( .D(n6815), .CLK(clk), .Q(arr[57]) );
  DFFPOSX1 arr_reg_1__23_ ( .D(n6814), .CLK(clk), .Q(arr[56]) );
  DFFPOSX1 arr_reg_1__22_ ( .D(n6813), .CLK(clk), .Q(arr[55]) );
  DFFPOSX1 arr_reg_1__21_ ( .D(n6812), .CLK(clk), .Q(arr[54]) );
  DFFPOSX1 arr_reg_1__20_ ( .D(n6811), .CLK(clk), .Q(arr[53]) );
  DFFPOSX1 arr_reg_1__19_ ( .D(n6810), .CLK(clk), .Q(arr[52]) );
  DFFPOSX1 arr_reg_1__18_ ( .D(n6809), .CLK(clk), .Q(arr[51]) );
  DFFPOSX1 arr_reg_1__17_ ( .D(n6808), .CLK(clk), .Q(arr[50]) );
  DFFPOSX1 arr_reg_1__16_ ( .D(n6807), .CLK(clk), .Q(arr[49]) );
  DFFPOSX1 arr_reg_1__15_ ( .D(n6806), .CLK(clk), .Q(arr[48]) );
  DFFPOSX1 arr_reg_1__14_ ( .D(n6805), .CLK(clk), .Q(arr[47]) );
  DFFPOSX1 arr_reg_1__13_ ( .D(n6804), .CLK(clk), .Q(arr[46]) );
  DFFPOSX1 arr_reg_1__12_ ( .D(n6803), .CLK(clk), .Q(arr[45]) );
  DFFPOSX1 arr_reg_1__11_ ( .D(n6802), .CLK(clk), .Q(arr[44]) );
  DFFPOSX1 arr_reg_1__10_ ( .D(n6801), .CLK(clk), .Q(arr[43]) );
  DFFPOSX1 arr_reg_1__9_ ( .D(n6800), .CLK(clk), .Q(arr[42]) );
  DFFPOSX1 arr_reg_1__8_ ( .D(n6799), .CLK(clk), .Q(arr[41]) );
  DFFPOSX1 arr_reg_1__7_ ( .D(n6798), .CLK(clk), .Q(arr[40]) );
  DFFPOSX1 arr_reg_1__6_ ( .D(n6797), .CLK(clk), .Q(arr[39]) );
  DFFPOSX1 arr_reg_1__5_ ( .D(n6796), .CLK(clk), .Q(arr[38]) );
  DFFPOSX1 arr_reg_1__4_ ( .D(n6795), .CLK(clk), .Q(arr[37]) );
  DFFPOSX1 arr_reg_1__3_ ( .D(n6794), .CLK(clk), .Q(arr[36]) );
  DFFPOSX1 arr_reg_1__2_ ( .D(n6793), .CLK(clk), .Q(arr[35]) );
  DFFPOSX1 arr_reg_1__1_ ( .D(n6792), .CLK(clk), .Q(arr[34]) );
  DFFPOSX1 arr_reg_1__0_ ( .D(n6791), .CLK(clk), .Q(arr[33]) );
  DFFPOSX1 arr_reg_0__32_ ( .D(n6790), .CLK(clk), .Q(arr[32]) );
  DFFPOSX1 arr_reg_0__31_ ( .D(n6789), .CLK(clk), .Q(arr[31]) );
  DFFPOSX1 arr_reg_0__30_ ( .D(n6788), .CLK(clk), .Q(arr[30]) );
  DFFPOSX1 arr_reg_0__29_ ( .D(n6787), .CLK(clk), .Q(arr[29]) );
  DFFPOSX1 arr_reg_0__28_ ( .D(n6786), .CLK(clk), .Q(arr[28]) );
  DFFPOSX1 arr_reg_0__27_ ( .D(n6785), .CLK(clk), .Q(arr[27]) );
  DFFPOSX1 arr_reg_0__26_ ( .D(n6784), .CLK(clk), .Q(arr[26]) );
  DFFPOSX1 arr_reg_0__25_ ( .D(n6783), .CLK(clk), .Q(arr[25]) );
  DFFPOSX1 arr_reg_0__24_ ( .D(n6782), .CLK(clk), .Q(arr[24]) );
  DFFPOSX1 arr_reg_0__23_ ( .D(n6781), .CLK(clk), .Q(arr[23]) );
  DFFPOSX1 arr_reg_0__22_ ( .D(n6780), .CLK(clk), .Q(arr[22]) );
  DFFPOSX1 arr_reg_0__21_ ( .D(n6779), .CLK(clk), .Q(arr[21]) );
  DFFPOSX1 arr_reg_0__20_ ( .D(n6778), .CLK(clk), .Q(arr[20]) );
  DFFPOSX1 arr_reg_0__19_ ( .D(n6777), .CLK(clk), .Q(arr[19]) );
  DFFPOSX1 arr_reg_0__18_ ( .D(n6776), .CLK(clk), .Q(arr[18]) );
  DFFPOSX1 arr_reg_0__17_ ( .D(n6775), .CLK(clk), .Q(arr[17]) );
  DFFPOSX1 arr_reg_0__16_ ( .D(n6774), .CLK(clk), .Q(arr[16]) );
  DFFPOSX1 arr_reg_0__15_ ( .D(n6773), .CLK(clk), .Q(arr[15]) );
  DFFPOSX1 arr_reg_0__14_ ( .D(n6772), .CLK(clk), .Q(arr[14]) );
  DFFPOSX1 arr_reg_0__13_ ( .D(n6771), .CLK(clk), .Q(arr[13]) );
  DFFPOSX1 arr_reg_0__12_ ( .D(n6770), .CLK(clk), .Q(arr[12]) );
  DFFPOSX1 arr_reg_0__11_ ( .D(n6769), .CLK(clk), .Q(arr[11]) );
  DFFPOSX1 arr_reg_0__10_ ( .D(n6768), .CLK(clk), .Q(arr[10]) );
  DFFPOSX1 arr_reg_0__9_ ( .D(n6767), .CLK(clk), .Q(arr[9]) );
  DFFPOSX1 arr_reg_0__8_ ( .D(n6766), .CLK(clk), .Q(arr[8]) );
  DFFPOSX1 arr_reg_0__7_ ( .D(n6765), .CLK(clk), .Q(arr[7]) );
  DFFPOSX1 arr_reg_0__6_ ( .D(n6764), .CLK(clk), .Q(arr[6]) );
  DFFPOSX1 arr_reg_0__5_ ( .D(n6763), .CLK(clk), .Q(arr[5]) );
  DFFPOSX1 arr_reg_0__4_ ( .D(n6762), .CLK(clk), .Q(arr[4]) );
  DFFPOSX1 arr_reg_0__3_ ( .D(n6761), .CLK(clk), .Q(arr[3]) );
  DFFPOSX1 arr_reg_0__2_ ( .D(n6760), .CLK(clk), .Q(arr[2]) );
  DFFPOSX1 arr_reg_0__1_ ( .D(n6759), .CLK(clk), .Q(arr[1]) );
  DFFPOSX1 arr_reg_0__0_ ( .D(n6758), .CLK(clk), .Q(arr[0]) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n6757), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n6756), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n6755), .CLK(clk), .Q(n15) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n6754), .CLK(clk), .Q(n16) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n6753), .CLK(clk), .Q(n17) );
  DFFPOSX1 rd_ptr_reg_5_ ( .D(n6752), .CLK(clk), .Q(n18) );
  AOI22X1 U4 ( .A(n2218), .B(n4458), .C(n18), .D(n4459), .Y(n4457) );
  AOI22X1 U6 ( .A(n2217), .B(n4458), .C(n17), .D(n4459), .Y(n4460) );
  AOI22X1 U8 ( .A(n2216), .B(n4458), .C(n16), .D(n4459), .Y(n4461) );
  AOI22X1 U10 ( .A(n2215), .B(n4458), .C(n15), .D(n4459), .Y(n4462) );
  AOI22X1 U12 ( .A(n2214), .B(n4458), .C(n14), .D(n4459), .Y(n4463) );
  AOI22X1 U14 ( .A(n2213), .B(n4458), .C(n13), .D(n4459), .Y(n4464) );
  NOR2X1 U15 ( .A(n4459), .B(reset), .Y(n4458) );
  OAI21X1 U17 ( .A(n2814), .B(n4467), .C(n4468), .Y(n6758) );
  NAND2X1 U18 ( .A(arr[0]), .B(n2816), .Y(n4468) );
  OAI21X1 U19 ( .A(n2814), .B(n4469), .C(n4470), .Y(n6759) );
  NAND2X1 U20 ( .A(arr[1]), .B(n2816), .Y(n4470) );
  OAI21X1 U21 ( .A(n2814), .B(n4471), .C(n4472), .Y(n6760) );
  NAND2X1 U22 ( .A(arr[2]), .B(n2816), .Y(n4472) );
  OAI21X1 U23 ( .A(n2814), .B(n4473), .C(n4474), .Y(n6761) );
  NAND2X1 U24 ( .A(arr[3]), .B(n2816), .Y(n4474) );
  OAI21X1 U25 ( .A(n2815), .B(n4475), .C(n4476), .Y(n6762) );
  NAND2X1 U26 ( .A(arr[4]), .B(n2816), .Y(n4476) );
  OAI21X1 U27 ( .A(n2815), .B(n4477), .C(n4478), .Y(n6763) );
  NAND2X1 U28 ( .A(arr[5]), .B(n2816), .Y(n4478) );
  OAI21X1 U29 ( .A(n2815), .B(n4479), .C(n4480), .Y(n6764) );
  NAND2X1 U30 ( .A(arr[6]), .B(n2814), .Y(n4480) );
  OAI21X1 U31 ( .A(n2816), .B(n4481), .C(n4482), .Y(n6765) );
  NAND2X1 U32 ( .A(arr[7]), .B(n2816), .Y(n4482) );
  OAI21X1 U33 ( .A(n2815), .B(n4483), .C(n4484), .Y(n6766) );
  NAND2X1 U34 ( .A(arr[8]), .B(n2816), .Y(n4484) );
  OAI21X1 U35 ( .A(n2816), .B(n4485), .C(n4486), .Y(n6767) );
  NAND2X1 U36 ( .A(arr[9]), .B(n2815), .Y(n4486) );
  OAI21X1 U37 ( .A(n2816), .B(n4487), .C(n4488), .Y(n6768) );
  NAND2X1 U38 ( .A(arr[10]), .B(n2814), .Y(n4488) );
  OAI21X1 U39 ( .A(n2815), .B(n4489), .C(n4490), .Y(n6769) );
  NAND2X1 U40 ( .A(arr[11]), .B(n2815), .Y(n4490) );
  OAI21X1 U41 ( .A(n2816), .B(n4491), .C(n4492), .Y(n6770) );
  NAND2X1 U42 ( .A(arr[12]), .B(n2815), .Y(n4492) );
  OAI21X1 U43 ( .A(n2816), .B(n4493), .C(n4494), .Y(n6771) );
  NAND2X1 U44 ( .A(arr[13]), .B(n2814), .Y(n4494) );
  OAI21X1 U45 ( .A(n2815), .B(n4495), .C(n4496), .Y(n6772) );
  NAND2X1 U46 ( .A(arr[14]), .B(n2816), .Y(n4496) );
  OAI21X1 U47 ( .A(n2816), .B(n4497), .C(n4498), .Y(n6773) );
  NAND2X1 U48 ( .A(arr[15]), .B(n2816), .Y(n4498) );
  OAI21X1 U49 ( .A(n2816), .B(n4499), .C(n4500), .Y(n6774) );
  NAND2X1 U50 ( .A(arr[16]), .B(n2816), .Y(n4500) );
  OAI21X1 U51 ( .A(n2815), .B(n4501), .C(n4502), .Y(n6775) );
  NAND2X1 U52 ( .A(arr[17]), .B(n2814), .Y(n4502) );
  OAI21X1 U53 ( .A(n2815), .B(n4503), .C(n4504), .Y(n6776) );
  NAND2X1 U54 ( .A(arr[18]), .B(n2816), .Y(n4504) );
  OAI21X1 U55 ( .A(n2815), .B(n4505), .C(n4506), .Y(n6777) );
  NAND2X1 U56 ( .A(arr[19]), .B(n2814), .Y(n4506) );
  OAI21X1 U57 ( .A(n2815), .B(n4507), .C(n4508), .Y(n6778) );
  NAND2X1 U58 ( .A(arr[20]), .B(n2815), .Y(n4508) );
  OAI21X1 U59 ( .A(n2815), .B(n4509), .C(n4510), .Y(n6779) );
  NAND2X1 U60 ( .A(arr[21]), .B(n2816), .Y(n4510) );
  OAI21X1 U61 ( .A(n2815), .B(n4511), .C(n4512), .Y(n6780) );
  NAND2X1 U62 ( .A(arr[22]), .B(n2816), .Y(n4512) );
  OAI21X1 U63 ( .A(n2814), .B(n4513), .C(n4514), .Y(n6781) );
  NAND2X1 U64 ( .A(arr[23]), .B(n2816), .Y(n4514) );
  OAI21X1 U65 ( .A(n2815), .B(n4515), .C(n4516), .Y(n6782) );
  NAND2X1 U66 ( .A(arr[24]), .B(n2815), .Y(n4516) );
  OAI21X1 U67 ( .A(n2814), .B(n4517), .C(n4518), .Y(n6783) );
  NAND2X1 U68 ( .A(arr[25]), .B(n2814), .Y(n4518) );
  OAI21X1 U69 ( .A(n2814), .B(n4519), .C(n4520), .Y(n6784) );
  NAND2X1 U70 ( .A(arr[26]), .B(n2815), .Y(n4520) );
  OAI21X1 U71 ( .A(n2814), .B(n4521), .C(n4522), .Y(n6785) );
  NAND2X1 U72 ( .A(arr[27]), .B(n2816), .Y(n4522) );
  OAI21X1 U73 ( .A(n2814), .B(n4523), .C(n4524), .Y(n6786) );
  NAND2X1 U74 ( .A(arr[28]), .B(n2815), .Y(n4524) );
  OAI21X1 U75 ( .A(n2814), .B(n4525), .C(n4526), .Y(n6787) );
  NAND2X1 U76 ( .A(arr[29]), .B(n2814), .Y(n4526) );
  OAI21X1 U77 ( .A(n2814), .B(n4527), .C(n4528), .Y(n6788) );
  NAND2X1 U78 ( .A(arr[30]), .B(n2815), .Y(n4528) );
  OAI21X1 U79 ( .A(n2814), .B(n4529), .C(n4530), .Y(n6789) );
  NAND2X1 U80 ( .A(arr[31]), .B(n2816), .Y(n4530) );
  OAI21X1 U81 ( .A(n2814), .B(n4531), .C(n4532), .Y(n6790) );
  NAND2X1 U82 ( .A(arr[32]), .B(n2814), .Y(n4532) );
  OAI21X1 U84 ( .A(n4467), .B(n2813), .C(n4536), .Y(n6791) );
  NAND2X1 U85 ( .A(arr[33]), .B(n2812), .Y(n4536) );
  OAI21X1 U86 ( .A(n4469), .B(n2811), .C(n4537), .Y(n6792) );
  NAND2X1 U87 ( .A(arr[34]), .B(n2812), .Y(n4537) );
  OAI21X1 U88 ( .A(n4471), .B(n2811), .C(n4538), .Y(n6793) );
  NAND2X1 U89 ( .A(arr[35]), .B(n2812), .Y(n4538) );
  OAI21X1 U90 ( .A(n4473), .B(n2811), .C(n4539), .Y(n6794) );
  NAND2X1 U91 ( .A(arr[36]), .B(n2812), .Y(n4539) );
  OAI21X1 U92 ( .A(n4475), .B(n2811), .C(n4540), .Y(n6795) );
  NAND2X1 U93 ( .A(arr[37]), .B(n2812), .Y(n4540) );
  OAI21X1 U94 ( .A(n4477), .B(n2811), .C(n4541), .Y(n6796) );
  NAND2X1 U95 ( .A(arr[38]), .B(n2813), .Y(n4541) );
  OAI21X1 U96 ( .A(n4479), .B(n2811), .C(n4542), .Y(n6797) );
  NAND2X1 U97 ( .A(arr[39]), .B(n2813), .Y(n4542) );
  OAI21X1 U98 ( .A(n4481), .B(n2812), .C(n4543), .Y(n6798) );
  NAND2X1 U99 ( .A(arr[40]), .B(n2812), .Y(n4543) );
  OAI21X1 U100 ( .A(n4483), .B(n2811), .C(n4544), .Y(n6799) );
  NAND2X1 U101 ( .A(arr[41]), .B(n2812), .Y(n4544) );
  OAI21X1 U102 ( .A(n4485), .B(n2812), .C(n4545), .Y(n6800) );
  NAND2X1 U103 ( .A(arr[42]), .B(n2813), .Y(n4545) );
  OAI21X1 U104 ( .A(n4487), .B(n2812), .C(n4546), .Y(n6801) );
  NAND2X1 U105 ( .A(arr[43]), .B(n2813), .Y(n4546) );
  OAI21X1 U106 ( .A(n4489), .B(n2811), .C(n4547), .Y(n6802) );
  NAND2X1 U107 ( .A(arr[44]), .B(n2813), .Y(n4547) );
  OAI21X1 U108 ( .A(n4491), .B(n2812), .C(n4548), .Y(n6803) );
  NAND2X1 U109 ( .A(arr[45]), .B(n2813), .Y(n4548) );
  OAI21X1 U110 ( .A(n4493), .B(n2812), .C(n4549), .Y(n6804) );
  NAND2X1 U111 ( .A(arr[46]), .B(n2813), .Y(n4549) );
  OAI21X1 U112 ( .A(n4495), .B(n2811), .C(n4550), .Y(n6805) );
  NAND2X1 U113 ( .A(arr[47]), .B(n2813), .Y(n4550) );
  OAI21X1 U114 ( .A(n4497), .B(n2812), .C(n4551), .Y(n6806) );
  NAND2X1 U115 ( .A(arr[48]), .B(n2813), .Y(n4551) );
  OAI21X1 U116 ( .A(n4499), .B(n2812), .C(n4552), .Y(n6807) );
  NAND2X1 U117 ( .A(arr[49]), .B(n2813), .Y(n4552) );
  OAI21X1 U118 ( .A(n4501), .B(n2811), .C(n4553), .Y(n6808) );
  NAND2X1 U119 ( .A(arr[50]), .B(n2813), .Y(n4553) );
  OAI21X1 U120 ( .A(n4503), .B(n2811), .C(n4554), .Y(n6809) );
  NAND2X1 U121 ( .A(arr[51]), .B(n2813), .Y(n4554) );
  OAI21X1 U122 ( .A(n4505), .B(n2811), .C(n4555), .Y(n6810) );
  NAND2X1 U123 ( .A(arr[52]), .B(n2813), .Y(n4555) );
  OAI21X1 U124 ( .A(n4507), .B(n2811), .C(n4556), .Y(n6811) );
  NAND2X1 U125 ( .A(arr[53]), .B(n2813), .Y(n4556) );
  OAI21X1 U126 ( .A(n4509), .B(n2811), .C(n4557), .Y(n6812) );
  NAND2X1 U127 ( .A(arr[54]), .B(n2813), .Y(n4557) );
  OAI21X1 U128 ( .A(n4511), .B(n2811), .C(n4558), .Y(n6813) );
  NAND2X1 U129 ( .A(arr[55]), .B(n2813), .Y(n4558) );
  OAI21X1 U130 ( .A(n4513), .B(n2813), .C(n4559), .Y(n6814) );
  NAND2X1 U131 ( .A(arr[56]), .B(n2813), .Y(n4559) );
  OAI21X1 U132 ( .A(n4515), .B(n2811), .C(n4560), .Y(n6815) );
  NAND2X1 U133 ( .A(arr[57]), .B(n2813), .Y(n4560) );
  OAI21X1 U134 ( .A(n4517), .B(n2812), .C(n4561), .Y(n6816) );
  NAND2X1 U135 ( .A(arr[58]), .B(n2813), .Y(n4561) );
  OAI21X1 U136 ( .A(n4519), .B(n2811), .C(n4562), .Y(n6817) );
  NAND2X1 U137 ( .A(arr[59]), .B(n2812), .Y(n4562) );
  OAI21X1 U138 ( .A(n4521), .B(n2812), .C(n4563), .Y(n6818) );
  NAND2X1 U139 ( .A(arr[60]), .B(n2813), .Y(n4563) );
  OAI21X1 U140 ( .A(n4523), .B(n2811), .C(n4564), .Y(n6819) );
  NAND2X1 U141 ( .A(arr[61]), .B(n2812), .Y(n4564) );
  OAI21X1 U142 ( .A(n4525), .B(n2811), .C(n4565), .Y(n6820) );
  NAND2X1 U143 ( .A(arr[62]), .B(n2813), .Y(n4565) );
  OAI21X1 U144 ( .A(n4527), .B(n2811), .C(n4566), .Y(n6821) );
  NAND2X1 U145 ( .A(arr[63]), .B(n2812), .Y(n4566) );
  OAI21X1 U146 ( .A(n4529), .B(n2811), .C(n4567), .Y(n6822) );
  NAND2X1 U147 ( .A(arr[64]), .B(n2812), .Y(n4567) );
  OAI21X1 U148 ( .A(n4531), .B(n2811), .C(n4568), .Y(n6823) );
  NAND2X1 U149 ( .A(arr[65]), .B(n2813), .Y(n4568) );
  OAI21X1 U151 ( .A(n4467), .B(n2808), .C(n4571), .Y(n6824) );
  NAND2X1 U152 ( .A(arr[66]), .B(n2810), .Y(n4571) );
  OAI21X1 U153 ( .A(n4469), .B(n2808), .C(n4572), .Y(n6825) );
  NAND2X1 U154 ( .A(arr[67]), .B(n2810), .Y(n4572) );
  OAI21X1 U155 ( .A(n4471), .B(n2808), .C(n4573), .Y(n6826) );
  NAND2X1 U156 ( .A(arr[68]), .B(n2810), .Y(n4573) );
  OAI21X1 U157 ( .A(n4473), .B(n2808), .C(n4574), .Y(n6827) );
  NAND2X1 U158 ( .A(arr[69]), .B(n2810), .Y(n4574) );
  OAI21X1 U159 ( .A(n4475), .B(n2809), .C(n4575), .Y(n6828) );
  NAND2X1 U160 ( .A(arr[70]), .B(n2810), .Y(n4575) );
  OAI21X1 U161 ( .A(n4477), .B(n2809), .C(n4576), .Y(n6829) );
  NAND2X1 U162 ( .A(arr[71]), .B(n2809), .Y(n4576) );
  OAI21X1 U163 ( .A(n4479), .B(n2809), .C(n4577), .Y(n6830) );
  NAND2X1 U164 ( .A(arr[72]), .B(n2810), .Y(n4577) );
  OAI21X1 U165 ( .A(n4481), .B(n2810), .C(n4578), .Y(n6831) );
  NAND2X1 U166 ( .A(arr[73]), .B(n2810), .Y(n4578) );
  OAI21X1 U167 ( .A(n4483), .B(n2809), .C(n4579), .Y(n6832) );
  NAND2X1 U168 ( .A(arr[74]), .B(n2810), .Y(n4579) );
  OAI21X1 U169 ( .A(n4485), .B(n2810), .C(n4580), .Y(n6833) );
  NAND2X1 U170 ( .A(arr[75]), .B(n2808), .Y(n4580) );
  OAI21X1 U171 ( .A(n4487), .B(n2810), .C(n4581), .Y(n6834) );
  NAND2X1 U172 ( .A(arr[76]), .B(n2810), .Y(n4581) );
  OAI21X1 U173 ( .A(n4489), .B(n2809), .C(n4582), .Y(n6835) );
  NAND2X1 U174 ( .A(arr[77]), .B(n2808), .Y(n4582) );
  OAI21X1 U175 ( .A(n4491), .B(n2810), .C(n4583), .Y(n6836) );
  NAND2X1 U176 ( .A(arr[78]), .B(n2809), .Y(n4583) );
  OAI21X1 U177 ( .A(n4493), .B(n2810), .C(n4584), .Y(n6837) );
  NAND2X1 U178 ( .A(arr[79]), .B(n2809), .Y(n4584) );
  OAI21X1 U179 ( .A(n4495), .B(n2809), .C(n4585), .Y(n6838) );
  NAND2X1 U180 ( .A(arr[80]), .B(n2810), .Y(n4585) );
  OAI21X1 U181 ( .A(n4497), .B(n2810), .C(n4586), .Y(n6839) );
  NAND2X1 U182 ( .A(arr[81]), .B(n2808), .Y(n4586) );
  OAI21X1 U183 ( .A(n4499), .B(n2810), .C(n4587), .Y(n6840) );
  NAND2X1 U184 ( .A(arr[82]), .B(n2810), .Y(n4587) );
  OAI21X1 U185 ( .A(n4501), .B(n2809), .C(n4588), .Y(n6841) );
  NAND2X1 U186 ( .A(arr[83]), .B(n2808), .Y(n4588) );
  OAI21X1 U187 ( .A(n4503), .B(n2809), .C(n4589), .Y(n6842) );
  NAND2X1 U188 ( .A(arr[84]), .B(n2809), .Y(n4589) );
  OAI21X1 U189 ( .A(n4505), .B(n2809), .C(n4590), .Y(n6843) );
  NAND2X1 U190 ( .A(arr[85]), .B(n2810), .Y(n4590) );
  OAI21X1 U191 ( .A(n4507), .B(n2809), .C(n4591), .Y(n6844) );
  NAND2X1 U192 ( .A(arr[86]), .B(n2808), .Y(n4591) );
  OAI21X1 U193 ( .A(n4509), .B(n2809), .C(n4592), .Y(n6845) );
  NAND2X1 U194 ( .A(arr[87]), .B(n2809), .Y(n4592) );
  OAI21X1 U195 ( .A(n4511), .B(n2809), .C(n4593), .Y(n6846) );
  NAND2X1 U196 ( .A(arr[88]), .B(n2810), .Y(n4593) );
  OAI21X1 U197 ( .A(n4513), .B(n2808), .C(n4594), .Y(n6847) );
  NAND2X1 U198 ( .A(arr[89]), .B(n2810), .Y(n4594) );
  OAI21X1 U199 ( .A(n4515), .B(n2809), .C(n4595), .Y(n6848) );
  NAND2X1 U200 ( .A(arr[90]), .B(n2810), .Y(n4595) );
  OAI21X1 U201 ( .A(n4517), .B(n2808), .C(n4596), .Y(n6849) );
  NAND2X1 U202 ( .A(arr[91]), .B(n2809), .Y(n4596) );
  OAI21X1 U203 ( .A(n4519), .B(n2808), .C(n4597), .Y(n6850) );
  NAND2X1 U204 ( .A(arr[92]), .B(n2808), .Y(n4597) );
  OAI21X1 U205 ( .A(n4521), .B(n2808), .C(n4598), .Y(n6851) );
  NAND2X1 U206 ( .A(arr[93]), .B(n2810), .Y(n4598) );
  OAI21X1 U207 ( .A(n4523), .B(n2808), .C(n4599), .Y(n6852) );
  NAND2X1 U208 ( .A(arr[94]), .B(n2809), .Y(n4599) );
  OAI21X1 U209 ( .A(n4525), .B(n2808), .C(n4600), .Y(n6853) );
  NAND2X1 U210 ( .A(arr[95]), .B(n2809), .Y(n4600) );
  OAI21X1 U211 ( .A(n4527), .B(n2808), .C(n4601), .Y(n6854) );
  NAND2X1 U212 ( .A(arr[96]), .B(n2808), .Y(n4601) );
  OAI21X1 U213 ( .A(n4529), .B(n2808), .C(n4602), .Y(n6855) );
  NAND2X1 U214 ( .A(arr[97]), .B(n2810), .Y(n4602) );
  OAI21X1 U215 ( .A(n4531), .B(n2808), .C(n4603), .Y(n6856) );
  NAND2X1 U216 ( .A(arr[98]), .B(n2808), .Y(n4603) );
  OAI21X1 U218 ( .A(n4467), .B(n2807), .C(n4606), .Y(n6857) );
  NAND2X1 U219 ( .A(arr[99]), .B(n2806), .Y(n4606) );
  OAI21X1 U220 ( .A(n4469), .B(n2805), .C(n4607), .Y(n6858) );
  NAND2X1 U221 ( .A(arr[100]), .B(n2806), .Y(n4607) );
  OAI21X1 U222 ( .A(n4471), .B(n2805), .C(n4608), .Y(n6859) );
  NAND2X1 U223 ( .A(arr[101]), .B(n2806), .Y(n4608) );
  OAI21X1 U224 ( .A(n4473), .B(n2805), .C(n4609), .Y(n6860) );
  NAND2X1 U225 ( .A(arr[102]), .B(n2806), .Y(n4609) );
  OAI21X1 U226 ( .A(n4475), .B(n2805), .C(n4610), .Y(n6861) );
  NAND2X1 U227 ( .A(arr[103]), .B(n2806), .Y(n4610) );
  OAI21X1 U228 ( .A(n4477), .B(n2805), .C(n4611), .Y(n6862) );
  NAND2X1 U229 ( .A(arr[104]), .B(n2807), .Y(n4611) );
  OAI21X1 U230 ( .A(n4479), .B(n2805), .C(n4612), .Y(n6863) );
  NAND2X1 U231 ( .A(arr[105]), .B(n2807), .Y(n4612) );
  OAI21X1 U232 ( .A(n4481), .B(n2806), .C(n4613), .Y(n6864) );
  NAND2X1 U233 ( .A(arr[106]), .B(n2806), .Y(n4613) );
  OAI21X1 U234 ( .A(n4483), .B(n2805), .C(n4614), .Y(n6865) );
  NAND2X1 U235 ( .A(arr[107]), .B(n2806), .Y(n4614) );
  OAI21X1 U236 ( .A(n4485), .B(n2806), .C(n4615), .Y(n6866) );
  NAND2X1 U237 ( .A(arr[108]), .B(n2807), .Y(n4615) );
  OAI21X1 U238 ( .A(n4487), .B(n2806), .C(n4616), .Y(n6867) );
  NAND2X1 U239 ( .A(arr[109]), .B(n2807), .Y(n4616) );
  OAI21X1 U240 ( .A(n4489), .B(n2805), .C(n4617), .Y(n6868) );
  NAND2X1 U241 ( .A(arr[110]), .B(n2807), .Y(n4617) );
  OAI21X1 U242 ( .A(n4491), .B(n2806), .C(n4618), .Y(n6869) );
  NAND2X1 U243 ( .A(arr[111]), .B(n2807), .Y(n4618) );
  OAI21X1 U244 ( .A(n4493), .B(n2806), .C(n4619), .Y(n6870) );
  NAND2X1 U245 ( .A(arr[112]), .B(n2807), .Y(n4619) );
  OAI21X1 U246 ( .A(n4495), .B(n2805), .C(n4620), .Y(n6871) );
  NAND2X1 U247 ( .A(arr[113]), .B(n2807), .Y(n4620) );
  OAI21X1 U248 ( .A(n4497), .B(n2806), .C(n4621), .Y(n6872) );
  NAND2X1 U249 ( .A(arr[114]), .B(n2807), .Y(n4621) );
  OAI21X1 U250 ( .A(n4499), .B(n2806), .C(n4622), .Y(n6873) );
  NAND2X1 U251 ( .A(arr[115]), .B(n2807), .Y(n4622) );
  OAI21X1 U252 ( .A(n4501), .B(n2805), .C(n4623), .Y(n6874) );
  NAND2X1 U253 ( .A(arr[116]), .B(n2807), .Y(n4623) );
  OAI21X1 U254 ( .A(n4503), .B(n2805), .C(n4624), .Y(n6875) );
  NAND2X1 U255 ( .A(arr[117]), .B(n2807), .Y(n4624) );
  OAI21X1 U256 ( .A(n4505), .B(n2805), .C(n4625), .Y(n6876) );
  NAND2X1 U257 ( .A(arr[118]), .B(n2807), .Y(n4625) );
  OAI21X1 U258 ( .A(n4507), .B(n2805), .C(n4626), .Y(n6877) );
  NAND2X1 U259 ( .A(arr[119]), .B(n2807), .Y(n4626) );
  OAI21X1 U260 ( .A(n4509), .B(n2805), .C(n4627), .Y(n6878) );
  NAND2X1 U261 ( .A(arr[120]), .B(n2807), .Y(n4627) );
  OAI21X1 U262 ( .A(n4511), .B(n2805), .C(n4628), .Y(n6879) );
  NAND2X1 U263 ( .A(arr[121]), .B(n2807), .Y(n4628) );
  OAI21X1 U264 ( .A(n4513), .B(n2807), .C(n4629), .Y(n6880) );
  NAND2X1 U265 ( .A(arr[122]), .B(n2807), .Y(n4629) );
  OAI21X1 U266 ( .A(n4515), .B(n2805), .C(n4630), .Y(n6881) );
  NAND2X1 U267 ( .A(arr[123]), .B(n2807), .Y(n4630) );
  OAI21X1 U268 ( .A(n4517), .B(n2806), .C(n4631), .Y(n6882) );
  NAND2X1 U269 ( .A(arr[124]), .B(n2807), .Y(n4631) );
  OAI21X1 U270 ( .A(n4519), .B(n2805), .C(n4632), .Y(n6883) );
  NAND2X1 U271 ( .A(arr[125]), .B(n2806), .Y(n4632) );
  OAI21X1 U272 ( .A(n4521), .B(n2806), .C(n4633), .Y(n6884) );
  NAND2X1 U273 ( .A(arr[126]), .B(n2807), .Y(n4633) );
  OAI21X1 U274 ( .A(n4523), .B(n2805), .C(n4634), .Y(n6885) );
  NAND2X1 U275 ( .A(arr[127]), .B(n2806), .Y(n4634) );
  OAI21X1 U276 ( .A(n4525), .B(n2805), .C(n4635), .Y(n6886) );
  NAND2X1 U277 ( .A(arr[128]), .B(n2807), .Y(n4635) );
  OAI21X1 U278 ( .A(n4527), .B(n2805), .C(n4636), .Y(n6887) );
  NAND2X1 U279 ( .A(arr[129]), .B(n2806), .Y(n4636) );
  OAI21X1 U280 ( .A(n4529), .B(n2805), .C(n4637), .Y(n6888) );
  NAND2X1 U281 ( .A(arr[130]), .B(n2806), .Y(n4637) );
  OAI21X1 U282 ( .A(n4531), .B(n2805), .C(n4638), .Y(n6889) );
  NAND2X1 U283 ( .A(arr[131]), .B(n2807), .Y(n4638) );
  OAI21X1 U285 ( .A(n4467), .B(n2802), .C(n4640), .Y(n6890) );
  NAND2X1 U286 ( .A(arr[132]), .B(n2804), .Y(n4640) );
  OAI21X1 U287 ( .A(n4469), .B(n2802), .C(n4641), .Y(n6891) );
  NAND2X1 U288 ( .A(arr[133]), .B(n2804), .Y(n4641) );
  OAI21X1 U289 ( .A(n4471), .B(n2802), .C(n4642), .Y(n6892) );
  NAND2X1 U290 ( .A(arr[134]), .B(n2804), .Y(n4642) );
  OAI21X1 U291 ( .A(n4473), .B(n2802), .C(n4643), .Y(n6893) );
  NAND2X1 U292 ( .A(arr[135]), .B(n2804), .Y(n4643) );
  OAI21X1 U293 ( .A(n4475), .B(n2803), .C(n4644), .Y(n6894) );
  NAND2X1 U294 ( .A(arr[136]), .B(n2804), .Y(n4644) );
  OAI21X1 U295 ( .A(n4477), .B(n2803), .C(n4645), .Y(n6895) );
  NAND2X1 U296 ( .A(arr[137]), .B(n2803), .Y(n4645) );
  OAI21X1 U297 ( .A(n4479), .B(n2803), .C(n4646), .Y(n6896) );
  NAND2X1 U298 ( .A(arr[138]), .B(n2804), .Y(n4646) );
  OAI21X1 U299 ( .A(n4481), .B(n2804), .C(n4647), .Y(n6897) );
  NAND2X1 U300 ( .A(arr[139]), .B(n2804), .Y(n4647) );
  OAI21X1 U301 ( .A(n4483), .B(n2803), .C(n4648), .Y(n6898) );
  NAND2X1 U302 ( .A(arr[140]), .B(n2804), .Y(n4648) );
  OAI21X1 U303 ( .A(n4485), .B(n2804), .C(n4649), .Y(n6899) );
  NAND2X1 U304 ( .A(arr[141]), .B(n2802), .Y(n4649) );
  OAI21X1 U305 ( .A(n4487), .B(n2804), .C(n4650), .Y(n6900) );
  NAND2X1 U306 ( .A(arr[142]), .B(n2804), .Y(n4650) );
  OAI21X1 U307 ( .A(n4489), .B(n2803), .C(n4651), .Y(n6901) );
  NAND2X1 U308 ( .A(arr[143]), .B(n2802), .Y(n4651) );
  OAI21X1 U309 ( .A(n4491), .B(n2804), .C(n4652), .Y(n6902) );
  NAND2X1 U310 ( .A(arr[144]), .B(n2803), .Y(n4652) );
  OAI21X1 U311 ( .A(n4493), .B(n2804), .C(n4653), .Y(n6903) );
  NAND2X1 U312 ( .A(arr[145]), .B(n2803), .Y(n4653) );
  OAI21X1 U313 ( .A(n4495), .B(n2803), .C(n4654), .Y(n6904) );
  NAND2X1 U314 ( .A(arr[146]), .B(n2804), .Y(n4654) );
  OAI21X1 U315 ( .A(n4497), .B(n2804), .C(n4655), .Y(n6905) );
  NAND2X1 U316 ( .A(arr[147]), .B(n2802), .Y(n4655) );
  OAI21X1 U317 ( .A(n4499), .B(n2804), .C(n4656), .Y(n6906) );
  NAND2X1 U318 ( .A(arr[148]), .B(n2804), .Y(n4656) );
  OAI21X1 U319 ( .A(n4501), .B(n2803), .C(n4657), .Y(n6907) );
  NAND2X1 U320 ( .A(arr[149]), .B(n2802), .Y(n4657) );
  OAI21X1 U321 ( .A(n4503), .B(n2803), .C(n4658), .Y(n6908) );
  NAND2X1 U322 ( .A(arr[150]), .B(n2803), .Y(n4658) );
  OAI21X1 U323 ( .A(n4505), .B(n2803), .C(n4659), .Y(n6909) );
  NAND2X1 U324 ( .A(arr[151]), .B(n2804), .Y(n4659) );
  OAI21X1 U325 ( .A(n4507), .B(n2803), .C(n4660), .Y(n6910) );
  NAND2X1 U326 ( .A(arr[152]), .B(n2802), .Y(n4660) );
  OAI21X1 U327 ( .A(n4509), .B(n2803), .C(n4661), .Y(n6911) );
  NAND2X1 U328 ( .A(arr[153]), .B(n2803), .Y(n4661) );
  OAI21X1 U329 ( .A(n4511), .B(n2803), .C(n4662), .Y(n6912) );
  NAND2X1 U330 ( .A(arr[154]), .B(n2804), .Y(n4662) );
  OAI21X1 U331 ( .A(n4513), .B(n2802), .C(n4663), .Y(n6913) );
  NAND2X1 U332 ( .A(arr[155]), .B(n2804), .Y(n4663) );
  OAI21X1 U333 ( .A(n4515), .B(n2803), .C(n4664), .Y(n6914) );
  NAND2X1 U334 ( .A(arr[156]), .B(n2804), .Y(n4664) );
  OAI21X1 U335 ( .A(n4517), .B(n2802), .C(n4665), .Y(n6915) );
  NAND2X1 U336 ( .A(arr[157]), .B(n2803), .Y(n4665) );
  OAI21X1 U337 ( .A(n4519), .B(n2802), .C(n4666), .Y(n6916) );
  NAND2X1 U338 ( .A(arr[158]), .B(n2802), .Y(n4666) );
  OAI21X1 U339 ( .A(n4521), .B(n2802), .C(n4667), .Y(n6917) );
  NAND2X1 U340 ( .A(arr[159]), .B(n2804), .Y(n4667) );
  OAI21X1 U341 ( .A(n4523), .B(n2802), .C(n4668), .Y(n6918) );
  NAND2X1 U342 ( .A(arr[160]), .B(n2803), .Y(n4668) );
  OAI21X1 U343 ( .A(n4525), .B(n2802), .C(n4669), .Y(n6919) );
  NAND2X1 U344 ( .A(arr[161]), .B(n2803), .Y(n4669) );
  OAI21X1 U345 ( .A(n4527), .B(n2802), .C(n4670), .Y(n6920) );
  NAND2X1 U346 ( .A(arr[162]), .B(n2802), .Y(n4670) );
  OAI21X1 U347 ( .A(n4529), .B(n2802), .C(n4671), .Y(n6921) );
  NAND2X1 U348 ( .A(arr[163]), .B(n2804), .Y(n4671) );
  OAI21X1 U349 ( .A(n4531), .B(n2802), .C(n4672), .Y(n6922) );
  NAND2X1 U350 ( .A(arr[164]), .B(n2802), .Y(n4672) );
  OAI21X1 U352 ( .A(n4467), .B(n2801), .C(n4675), .Y(n6923) );
  NAND2X1 U353 ( .A(arr[165]), .B(n2800), .Y(n4675) );
  OAI21X1 U354 ( .A(n4469), .B(n2799), .C(n4676), .Y(n6924) );
  NAND2X1 U355 ( .A(arr[166]), .B(n2800), .Y(n4676) );
  OAI21X1 U356 ( .A(n4471), .B(n2799), .C(n4677), .Y(n6925) );
  NAND2X1 U357 ( .A(arr[167]), .B(n2800), .Y(n4677) );
  OAI21X1 U358 ( .A(n4473), .B(n2799), .C(n4678), .Y(n6926) );
  NAND2X1 U359 ( .A(arr[168]), .B(n2800), .Y(n4678) );
  OAI21X1 U360 ( .A(n4475), .B(n2799), .C(n4679), .Y(n6927) );
  NAND2X1 U361 ( .A(arr[169]), .B(n2800), .Y(n4679) );
  OAI21X1 U362 ( .A(n4477), .B(n2799), .C(n4680), .Y(n6928) );
  NAND2X1 U363 ( .A(arr[170]), .B(n2801), .Y(n4680) );
  OAI21X1 U364 ( .A(n4479), .B(n2799), .C(n4681), .Y(n6929) );
  NAND2X1 U365 ( .A(arr[171]), .B(n2801), .Y(n4681) );
  OAI21X1 U366 ( .A(n4481), .B(n2800), .C(n4682), .Y(n6930) );
  NAND2X1 U367 ( .A(arr[172]), .B(n2800), .Y(n4682) );
  OAI21X1 U368 ( .A(n4483), .B(n2799), .C(n4683), .Y(n6931) );
  NAND2X1 U369 ( .A(arr[173]), .B(n2800), .Y(n4683) );
  OAI21X1 U370 ( .A(n4485), .B(n2800), .C(n4684), .Y(n6932) );
  NAND2X1 U371 ( .A(arr[174]), .B(n2801), .Y(n4684) );
  OAI21X1 U372 ( .A(n4487), .B(n2800), .C(n4685), .Y(n6933) );
  NAND2X1 U373 ( .A(arr[175]), .B(n2801), .Y(n4685) );
  OAI21X1 U374 ( .A(n4489), .B(n2799), .C(n4686), .Y(n6934) );
  NAND2X1 U375 ( .A(arr[176]), .B(n2801), .Y(n4686) );
  OAI21X1 U376 ( .A(n4491), .B(n2800), .C(n4687), .Y(n6935) );
  NAND2X1 U377 ( .A(arr[177]), .B(n2801), .Y(n4687) );
  OAI21X1 U378 ( .A(n4493), .B(n2800), .C(n4688), .Y(n6936) );
  NAND2X1 U379 ( .A(arr[178]), .B(n2801), .Y(n4688) );
  OAI21X1 U380 ( .A(n4495), .B(n2799), .C(n4689), .Y(n6937) );
  NAND2X1 U381 ( .A(arr[179]), .B(n2801), .Y(n4689) );
  OAI21X1 U382 ( .A(n4497), .B(n2800), .C(n4690), .Y(n6938) );
  NAND2X1 U383 ( .A(arr[180]), .B(n2801), .Y(n4690) );
  OAI21X1 U384 ( .A(n4499), .B(n2800), .C(n4691), .Y(n6939) );
  NAND2X1 U385 ( .A(arr[181]), .B(n2801), .Y(n4691) );
  OAI21X1 U386 ( .A(n4501), .B(n2799), .C(n4692), .Y(n6940) );
  NAND2X1 U387 ( .A(arr[182]), .B(n2801), .Y(n4692) );
  OAI21X1 U388 ( .A(n4503), .B(n2799), .C(n4693), .Y(n6941) );
  NAND2X1 U389 ( .A(arr[183]), .B(n2801), .Y(n4693) );
  OAI21X1 U390 ( .A(n4505), .B(n2799), .C(n4694), .Y(n6942) );
  NAND2X1 U391 ( .A(arr[184]), .B(n2801), .Y(n4694) );
  OAI21X1 U392 ( .A(n4507), .B(n2799), .C(n4695), .Y(n6943) );
  NAND2X1 U393 ( .A(arr[185]), .B(n2801), .Y(n4695) );
  OAI21X1 U394 ( .A(n4509), .B(n2799), .C(n4696), .Y(n6944) );
  NAND2X1 U395 ( .A(arr[186]), .B(n2801), .Y(n4696) );
  OAI21X1 U396 ( .A(n4511), .B(n2799), .C(n4697), .Y(n6945) );
  NAND2X1 U397 ( .A(arr[187]), .B(n2801), .Y(n4697) );
  OAI21X1 U398 ( .A(n4513), .B(n2801), .C(n4698), .Y(n6946) );
  NAND2X1 U399 ( .A(arr[188]), .B(n2801), .Y(n4698) );
  OAI21X1 U400 ( .A(n4515), .B(n2799), .C(n4699), .Y(n6947) );
  NAND2X1 U401 ( .A(arr[189]), .B(n2801), .Y(n4699) );
  OAI21X1 U402 ( .A(n4517), .B(n2800), .C(n4700), .Y(n6948) );
  NAND2X1 U403 ( .A(arr[190]), .B(n2801), .Y(n4700) );
  OAI21X1 U404 ( .A(n4519), .B(n2799), .C(n4701), .Y(n6949) );
  NAND2X1 U405 ( .A(arr[191]), .B(n2800), .Y(n4701) );
  OAI21X1 U406 ( .A(n4521), .B(n2800), .C(n4702), .Y(n6950) );
  NAND2X1 U407 ( .A(arr[192]), .B(n2801), .Y(n4702) );
  OAI21X1 U408 ( .A(n4523), .B(n2799), .C(n4703), .Y(n6951) );
  NAND2X1 U409 ( .A(arr[193]), .B(n2800), .Y(n4703) );
  OAI21X1 U410 ( .A(n4525), .B(n2799), .C(n4704), .Y(n6952) );
  NAND2X1 U411 ( .A(arr[194]), .B(n2801), .Y(n4704) );
  OAI21X1 U412 ( .A(n4527), .B(n2799), .C(n4705), .Y(n6953) );
  NAND2X1 U413 ( .A(arr[195]), .B(n2800), .Y(n4705) );
  OAI21X1 U414 ( .A(n4529), .B(n2799), .C(n4706), .Y(n6954) );
  NAND2X1 U415 ( .A(arr[196]), .B(n2800), .Y(n4706) );
  OAI21X1 U416 ( .A(n4531), .B(n2799), .C(n4707), .Y(n6955) );
  NAND2X1 U417 ( .A(arr[197]), .B(n2801), .Y(n4707) );
  OAI21X1 U419 ( .A(n4467), .B(n2796), .C(n4709), .Y(n6956) );
  NAND2X1 U420 ( .A(arr[198]), .B(n2798), .Y(n4709) );
  OAI21X1 U421 ( .A(n4469), .B(n2796), .C(n4710), .Y(n6957) );
  NAND2X1 U422 ( .A(arr[199]), .B(n2798), .Y(n4710) );
  OAI21X1 U423 ( .A(n4471), .B(n2796), .C(n4711), .Y(n6958) );
  NAND2X1 U424 ( .A(arr[200]), .B(n2798), .Y(n4711) );
  OAI21X1 U425 ( .A(n4473), .B(n2796), .C(n4712), .Y(n6959) );
  NAND2X1 U426 ( .A(arr[201]), .B(n2798), .Y(n4712) );
  OAI21X1 U427 ( .A(n4475), .B(n2797), .C(n4713), .Y(n6960) );
  NAND2X1 U428 ( .A(arr[202]), .B(n2798), .Y(n4713) );
  OAI21X1 U429 ( .A(n4477), .B(n2797), .C(n4714), .Y(n6961) );
  NAND2X1 U430 ( .A(arr[203]), .B(n2797), .Y(n4714) );
  OAI21X1 U431 ( .A(n4479), .B(n2797), .C(n4715), .Y(n6962) );
  NAND2X1 U432 ( .A(arr[204]), .B(n2798), .Y(n4715) );
  OAI21X1 U433 ( .A(n4481), .B(n2798), .C(n4716), .Y(n6963) );
  NAND2X1 U434 ( .A(arr[205]), .B(n2798), .Y(n4716) );
  OAI21X1 U435 ( .A(n4483), .B(n2797), .C(n4717), .Y(n6964) );
  NAND2X1 U436 ( .A(arr[206]), .B(n2798), .Y(n4717) );
  OAI21X1 U437 ( .A(n4485), .B(n2798), .C(n4718), .Y(n6965) );
  NAND2X1 U438 ( .A(arr[207]), .B(n2796), .Y(n4718) );
  OAI21X1 U439 ( .A(n4487), .B(n2798), .C(n4719), .Y(n6966) );
  NAND2X1 U440 ( .A(arr[208]), .B(n2798), .Y(n4719) );
  OAI21X1 U441 ( .A(n4489), .B(n2797), .C(n4720), .Y(n6967) );
  NAND2X1 U442 ( .A(arr[209]), .B(n2796), .Y(n4720) );
  OAI21X1 U443 ( .A(n4491), .B(n2798), .C(n4721), .Y(n6968) );
  NAND2X1 U444 ( .A(arr[210]), .B(n2797), .Y(n4721) );
  OAI21X1 U445 ( .A(n4493), .B(n2798), .C(n4722), .Y(n6969) );
  NAND2X1 U446 ( .A(arr[211]), .B(n2797), .Y(n4722) );
  OAI21X1 U447 ( .A(n4495), .B(n2797), .C(n4723), .Y(n6970) );
  NAND2X1 U448 ( .A(arr[212]), .B(n2798), .Y(n4723) );
  OAI21X1 U449 ( .A(n4497), .B(n2798), .C(n4724), .Y(n6971) );
  NAND2X1 U450 ( .A(arr[213]), .B(n2796), .Y(n4724) );
  OAI21X1 U451 ( .A(n4499), .B(n2798), .C(n4725), .Y(n6972) );
  NAND2X1 U452 ( .A(arr[214]), .B(n2798), .Y(n4725) );
  OAI21X1 U453 ( .A(n4501), .B(n2797), .C(n4726), .Y(n6973) );
  NAND2X1 U454 ( .A(arr[215]), .B(n2796), .Y(n4726) );
  OAI21X1 U455 ( .A(n4503), .B(n2797), .C(n4727), .Y(n6974) );
  NAND2X1 U456 ( .A(arr[216]), .B(n2797), .Y(n4727) );
  OAI21X1 U457 ( .A(n4505), .B(n2797), .C(n4728), .Y(n6975) );
  NAND2X1 U458 ( .A(arr[217]), .B(n2798), .Y(n4728) );
  OAI21X1 U459 ( .A(n4507), .B(n2797), .C(n4729), .Y(n6976) );
  NAND2X1 U460 ( .A(arr[218]), .B(n2796), .Y(n4729) );
  OAI21X1 U461 ( .A(n4509), .B(n2797), .C(n4730), .Y(n6977) );
  NAND2X1 U462 ( .A(arr[219]), .B(n2797), .Y(n4730) );
  OAI21X1 U463 ( .A(n4511), .B(n2797), .C(n4731), .Y(n6978) );
  NAND2X1 U464 ( .A(arr[220]), .B(n2798), .Y(n4731) );
  OAI21X1 U465 ( .A(n4513), .B(n2796), .C(n4732), .Y(n6979) );
  NAND2X1 U466 ( .A(arr[221]), .B(n2798), .Y(n4732) );
  OAI21X1 U467 ( .A(n4515), .B(n2797), .C(n4733), .Y(n6980) );
  NAND2X1 U468 ( .A(arr[222]), .B(n2798), .Y(n4733) );
  OAI21X1 U469 ( .A(n4517), .B(n2796), .C(n4734), .Y(n6981) );
  NAND2X1 U470 ( .A(arr[223]), .B(n2797), .Y(n4734) );
  OAI21X1 U471 ( .A(n4519), .B(n2796), .C(n4735), .Y(n6982) );
  NAND2X1 U472 ( .A(arr[224]), .B(n2796), .Y(n4735) );
  OAI21X1 U473 ( .A(n4521), .B(n2796), .C(n4736), .Y(n6983) );
  NAND2X1 U474 ( .A(arr[225]), .B(n2798), .Y(n4736) );
  OAI21X1 U475 ( .A(n4523), .B(n2796), .C(n4737), .Y(n6984) );
  NAND2X1 U476 ( .A(arr[226]), .B(n2797), .Y(n4737) );
  OAI21X1 U477 ( .A(n4525), .B(n2796), .C(n4738), .Y(n6985) );
  NAND2X1 U478 ( .A(arr[227]), .B(n2797), .Y(n4738) );
  OAI21X1 U479 ( .A(n4527), .B(n2796), .C(n4739), .Y(n6986) );
  NAND2X1 U480 ( .A(arr[228]), .B(n2796), .Y(n4739) );
  OAI21X1 U481 ( .A(n4529), .B(n2796), .C(n4740), .Y(n6987) );
  NAND2X1 U482 ( .A(arr[229]), .B(n2798), .Y(n4740) );
  OAI21X1 U483 ( .A(n4531), .B(n2796), .C(n4741), .Y(n6988) );
  NAND2X1 U484 ( .A(arr[230]), .B(n2796), .Y(n4741) );
  OAI21X1 U486 ( .A(n4467), .B(n2795), .C(n4744), .Y(n6989) );
  NAND2X1 U487 ( .A(arr[231]), .B(n2794), .Y(n4744) );
  OAI21X1 U488 ( .A(n4469), .B(n2793), .C(n4745), .Y(n6990) );
  NAND2X1 U489 ( .A(arr[232]), .B(n2794), .Y(n4745) );
  OAI21X1 U490 ( .A(n4471), .B(n2793), .C(n4746), .Y(n6991) );
  NAND2X1 U491 ( .A(arr[233]), .B(n2794), .Y(n4746) );
  OAI21X1 U492 ( .A(n4473), .B(n2793), .C(n4747), .Y(n6992) );
  NAND2X1 U493 ( .A(arr[234]), .B(n2794), .Y(n4747) );
  OAI21X1 U494 ( .A(n4475), .B(n2793), .C(n4748), .Y(n6993) );
  NAND2X1 U495 ( .A(arr[235]), .B(n2794), .Y(n4748) );
  OAI21X1 U496 ( .A(n4477), .B(n2793), .C(n4749), .Y(n6994) );
  NAND2X1 U497 ( .A(arr[236]), .B(n2795), .Y(n4749) );
  OAI21X1 U498 ( .A(n4479), .B(n2793), .C(n4750), .Y(n6995) );
  NAND2X1 U499 ( .A(arr[237]), .B(n2795), .Y(n4750) );
  OAI21X1 U500 ( .A(n4481), .B(n2794), .C(n4751), .Y(n6996) );
  NAND2X1 U501 ( .A(arr[238]), .B(n2794), .Y(n4751) );
  OAI21X1 U502 ( .A(n4483), .B(n2793), .C(n4752), .Y(n6997) );
  NAND2X1 U503 ( .A(arr[239]), .B(n2794), .Y(n4752) );
  OAI21X1 U504 ( .A(n4485), .B(n2794), .C(n4753), .Y(n6998) );
  NAND2X1 U505 ( .A(arr[240]), .B(n2795), .Y(n4753) );
  OAI21X1 U506 ( .A(n4487), .B(n2794), .C(n4754), .Y(n6999) );
  NAND2X1 U507 ( .A(arr[241]), .B(n2795), .Y(n4754) );
  OAI21X1 U508 ( .A(n4489), .B(n2793), .C(n4755), .Y(n7000) );
  NAND2X1 U509 ( .A(arr[242]), .B(n2795), .Y(n4755) );
  OAI21X1 U510 ( .A(n4491), .B(n2794), .C(n4756), .Y(n7001) );
  NAND2X1 U511 ( .A(arr[243]), .B(n2795), .Y(n4756) );
  OAI21X1 U512 ( .A(n4493), .B(n2794), .C(n4757), .Y(n7002) );
  NAND2X1 U513 ( .A(arr[244]), .B(n2795), .Y(n4757) );
  OAI21X1 U514 ( .A(n4495), .B(n2793), .C(n4758), .Y(n7003) );
  NAND2X1 U515 ( .A(arr[245]), .B(n2795), .Y(n4758) );
  OAI21X1 U516 ( .A(n4497), .B(n2794), .C(n4759), .Y(n7004) );
  NAND2X1 U517 ( .A(arr[246]), .B(n2795), .Y(n4759) );
  OAI21X1 U518 ( .A(n4499), .B(n2794), .C(n4760), .Y(n7005) );
  NAND2X1 U519 ( .A(arr[247]), .B(n2795), .Y(n4760) );
  OAI21X1 U520 ( .A(n4501), .B(n2793), .C(n4761), .Y(n7006) );
  NAND2X1 U521 ( .A(arr[248]), .B(n2795), .Y(n4761) );
  OAI21X1 U522 ( .A(n4503), .B(n2793), .C(n4762), .Y(n7007) );
  NAND2X1 U523 ( .A(arr[249]), .B(n2795), .Y(n4762) );
  OAI21X1 U524 ( .A(n4505), .B(n2793), .C(n4763), .Y(n7008) );
  NAND2X1 U525 ( .A(arr[250]), .B(n2795), .Y(n4763) );
  OAI21X1 U526 ( .A(n4507), .B(n2793), .C(n4764), .Y(n7009) );
  NAND2X1 U527 ( .A(arr[251]), .B(n2795), .Y(n4764) );
  OAI21X1 U528 ( .A(n4509), .B(n2793), .C(n4765), .Y(n7010) );
  NAND2X1 U529 ( .A(arr[252]), .B(n2795), .Y(n4765) );
  OAI21X1 U530 ( .A(n4511), .B(n2793), .C(n4766), .Y(n7011) );
  NAND2X1 U531 ( .A(arr[253]), .B(n2795), .Y(n4766) );
  OAI21X1 U532 ( .A(n4513), .B(n2795), .C(n4767), .Y(n7012) );
  NAND2X1 U533 ( .A(arr[254]), .B(n2795), .Y(n4767) );
  OAI21X1 U534 ( .A(n4515), .B(n2793), .C(n4768), .Y(n7013) );
  NAND2X1 U535 ( .A(arr[255]), .B(n2795), .Y(n4768) );
  OAI21X1 U536 ( .A(n4517), .B(n2794), .C(n4769), .Y(n7014) );
  NAND2X1 U537 ( .A(arr[256]), .B(n2795), .Y(n4769) );
  OAI21X1 U538 ( .A(n4519), .B(n2793), .C(n4770), .Y(n7015) );
  NAND2X1 U539 ( .A(arr[257]), .B(n2794), .Y(n4770) );
  OAI21X1 U540 ( .A(n4521), .B(n2794), .C(n4771), .Y(n7016) );
  NAND2X1 U541 ( .A(arr[258]), .B(n2795), .Y(n4771) );
  OAI21X1 U542 ( .A(n4523), .B(n2793), .C(n4772), .Y(n7017) );
  NAND2X1 U543 ( .A(arr[259]), .B(n2794), .Y(n4772) );
  OAI21X1 U544 ( .A(n4525), .B(n2793), .C(n4773), .Y(n7018) );
  NAND2X1 U545 ( .A(arr[260]), .B(n2795), .Y(n4773) );
  OAI21X1 U546 ( .A(n4527), .B(n2793), .C(n4774), .Y(n7019) );
  NAND2X1 U547 ( .A(arr[261]), .B(n2794), .Y(n4774) );
  OAI21X1 U548 ( .A(n4529), .B(n2793), .C(n4775), .Y(n7020) );
  NAND2X1 U549 ( .A(arr[262]), .B(n2794), .Y(n4775) );
  OAI21X1 U550 ( .A(n4531), .B(n2793), .C(n4776), .Y(n7021) );
  NAND2X1 U551 ( .A(arr[263]), .B(n2795), .Y(n4776) );
  OAI21X1 U553 ( .A(n4467), .B(n2790), .C(n4778), .Y(n7022) );
  NAND2X1 U554 ( .A(arr[264]), .B(n2792), .Y(n4778) );
  OAI21X1 U555 ( .A(n4469), .B(n2790), .C(n4779), .Y(n7023) );
  NAND2X1 U556 ( .A(arr[265]), .B(n2792), .Y(n4779) );
  OAI21X1 U557 ( .A(n4471), .B(n2790), .C(n4780), .Y(n7024) );
  NAND2X1 U558 ( .A(arr[266]), .B(n2792), .Y(n4780) );
  OAI21X1 U559 ( .A(n4473), .B(n2790), .C(n4781), .Y(n7025) );
  NAND2X1 U560 ( .A(arr[267]), .B(n2792), .Y(n4781) );
  OAI21X1 U561 ( .A(n4475), .B(n2791), .C(n4782), .Y(n7026) );
  NAND2X1 U562 ( .A(arr[268]), .B(n2792), .Y(n4782) );
  OAI21X1 U563 ( .A(n4477), .B(n2791), .C(n4783), .Y(n7027) );
  NAND2X1 U564 ( .A(arr[269]), .B(n2791), .Y(n4783) );
  OAI21X1 U565 ( .A(n4479), .B(n2791), .C(n4784), .Y(n7028) );
  NAND2X1 U566 ( .A(arr[270]), .B(n2792), .Y(n4784) );
  OAI21X1 U567 ( .A(n4481), .B(n2792), .C(n4785), .Y(n7029) );
  NAND2X1 U568 ( .A(arr[271]), .B(n2792), .Y(n4785) );
  OAI21X1 U569 ( .A(n4483), .B(n2791), .C(n4786), .Y(n7030) );
  NAND2X1 U570 ( .A(arr[272]), .B(n2792), .Y(n4786) );
  OAI21X1 U571 ( .A(n4485), .B(n2792), .C(n4787), .Y(n7031) );
  NAND2X1 U572 ( .A(arr[273]), .B(n2790), .Y(n4787) );
  OAI21X1 U573 ( .A(n4487), .B(n2792), .C(n4788), .Y(n7032) );
  NAND2X1 U574 ( .A(arr[274]), .B(n2792), .Y(n4788) );
  OAI21X1 U575 ( .A(n4489), .B(n2791), .C(n4789), .Y(n7033) );
  NAND2X1 U576 ( .A(arr[275]), .B(n2790), .Y(n4789) );
  OAI21X1 U577 ( .A(n4491), .B(n2792), .C(n4790), .Y(n7034) );
  NAND2X1 U578 ( .A(arr[276]), .B(n2791), .Y(n4790) );
  OAI21X1 U579 ( .A(n4493), .B(n2792), .C(n4791), .Y(n7035) );
  NAND2X1 U580 ( .A(arr[277]), .B(n2791), .Y(n4791) );
  OAI21X1 U581 ( .A(n4495), .B(n2791), .C(n4792), .Y(n7036) );
  NAND2X1 U582 ( .A(arr[278]), .B(n2792), .Y(n4792) );
  OAI21X1 U583 ( .A(n4497), .B(n2792), .C(n4793), .Y(n7037) );
  NAND2X1 U584 ( .A(arr[279]), .B(n2790), .Y(n4793) );
  OAI21X1 U585 ( .A(n4499), .B(n2792), .C(n4794), .Y(n7038) );
  NAND2X1 U586 ( .A(arr[280]), .B(n2792), .Y(n4794) );
  OAI21X1 U587 ( .A(n4501), .B(n2791), .C(n4795), .Y(n7039) );
  NAND2X1 U588 ( .A(arr[281]), .B(n2790), .Y(n4795) );
  OAI21X1 U589 ( .A(n4503), .B(n2791), .C(n4796), .Y(n7040) );
  NAND2X1 U590 ( .A(arr[282]), .B(n2791), .Y(n4796) );
  OAI21X1 U591 ( .A(n4505), .B(n2791), .C(n4797), .Y(n7041) );
  NAND2X1 U592 ( .A(arr[283]), .B(n2792), .Y(n4797) );
  OAI21X1 U593 ( .A(n4507), .B(n2791), .C(n4798), .Y(n7042) );
  NAND2X1 U594 ( .A(arr[284]), .B(n2790), .Y(n4798) );
  OAI21X1 U595 ( .A(n4509), .B(n2791), .C(n4799), .Y(n7043) );
  NAND2X1 U596 ( .A(arr[285]), .B(n2791), .Y(n4799) );
  OAI21X1 U597 ( .A(n4511), .B(n2791), .C(n4800), .Y(n7044) );
  NAND2X1 U598 ( .A(arr[286]), .B(n2792), .Y(n4800) );
  OAI21X1 U599 ( .A(n4513), .B(n2790), .C(n4801), .Y(n7045) );
  NAND2X1 U600 ( .A(arr[287]), .B(n2792), .Y(n4801) );
  OAI21X1 U601 ( .A(n4515), .B(n2791), .C(n4802), .Y(n7046) );
  NAND2X1 U602 ( .A(arr[288]), .B(n2792), .Y(n4802) );
  OAI21X1 U603 ( .A(n4517), .B(n2790), .C(n4803), .Y(n7047) );
  NAND2X1 U604 ( .A(arr[289]), .B(n2791), .Y(n4803) );
  OAI21X1 U605 ( .A(n4519), .B(n2790), .C(n4804), .Y(n7048) );
  NAND2X1 U606 ( .A(arr[290]), .B(n2790), .Y(n4804) );
  OAI21X1 U607 ( .A(n4521), .B(n2790), .C(n4805), .Y(n7049) );
  NAND2X1 U608 ( .A(arr[291]), .B(n2792), .Y(n4805) );
  OAI21X1 U609 ( .A(n4523), .B(n2790), .C(n4806), .Y(n7050) );
  NAND2X1 U610 ( .A(arr[292]), .B(n2791), .Y(n4806) );
  OAI21X1 U611 ( .A(n4525), .B(n2790), .C(n4807), .Y(n7051) );
  NAND2X1 U612 ( .A(arr[293]), .B(n2791), .Y(n4807) );
  OAI21X1 U613 ( .A(n4527), .B(n2790), .C(n4808), .Y(n7052) );
  NAND2X1 U614 ( .A(arr[294]), .B(n2790), .Y(n4808) );
  OAI21X1 U615 ( .A(n4529), .B(n2790), .C(n4809), .Y(n7053) );
  NAND2X1 U616 ( .A(arr[295]), .B(n2792), .Y(n4809) );
  OAI21X1 U617 ( .A(n4531), .B(n2790), .C(n4810), .Y(n7054) );
  NAND2X1 U618 ( .A(arr[296]), .B(n2790), .Y(n4810) );
  OAI21X1 U620 ( .A(n4467), .B(n2789), .C(n4813), .Y(n7055) );
  NAND2X1 U621 ( .A(arr[297]), .B(n2788), .Y(n4813) );
  OAI21X1 U622 ( .A(n4469), .B(n2787), .C(n4814), .Y(n7056) );
  NAND2X1 U623 ( .A(arr[298]), .B(n2788), .Y(n4814) );
  OAI21X1 U624 ( .A(n4471), .B(n2787), .C(n4815), .Y(n7057) );
  NAND2X1 U625 ( .A(arr[299]), .B(n2788), .Y(n4815) );
  OAI21X1 U626 ( .A(n4473), .B(n2787), .C(n4816), .Y(n7058) );
  NAND2X1 U627 ( .A(arr[300]), .B(n2788), .Y(n4816) );
  OAI21X1 U628 ( .A(n4475), .B(n2787), .C(n4817), .Y(n7059) );
  NAND2X1 U629 ( .A(arr[301]), .B(n2788), .Y(n4817) );
  OAI21X1 U630 ( .A(n4477), .B(n2787), .C(n4818), .Y(n7060) );
  NAND2X1 U631 ( .A(arr[302]), .B(n2789), .Y(n4818) );
  OAI21X1 U632 ( .A(n4479), .B(n2787), .C(n4819), .Y(n7061) );
  NAND2X1 U633 ( .A(arr[303]), .B(n2789), .Y(n4819) );
  OAI21X1 U634 ( .A(n4481), .B(n2788), .C(n4820), .Y(n7062) );
  NAND2X1 U635 ( .A(arr[304]), .B(n2788), .Y(n4820) );
  OAI21X1 U636 ( .A(n4483), .B(n2787), .C(n4821), .Y(n7063) );
  NAND2X1 U637 ( .A(arr[305]), .B(n2788), .Y(n4821) );
  OAI21X1 U638 ( .A(n4485), .B(n2788), .C(n4822), .Y(n7064) );
  NAND2X1 U639 ( .A(arr[306]), .B(n2789), .Y(n4822) );
  OAI21X1 U640 ( .A(n4487), .B(n2788), .C(n4823), .Y(n7065) );
  NAND2X1 U641 ( .A(arr[307]), .B(n2789), .Y(n4823) );
  OAI21X1 U642 ( .A(n4489), .B(n2787), .C(n4824), .Y(n7066) );
  NAND2X1 U643 ( .A(arr[308]), .B(n2789), .Y(n4824) );
  OAI21X1 U644 ( .A(n4491), .B(n2788), .C(n4825), .Y(n7067) );
  NAND2X1 U645 ( .A(arr[309]), .B(n2789), .Y(n4825) );
  OAI21X1 U646 ( .A(n4493), .B(n2788), .C(n4826), .Y(n7068) );
  NAND2X1 U647 ( .A(arr[310]), .B(n2789), .Y(n4826) );
  OAI21X1 U648 ( .A(n4495), .B(n2787), .C(n4827), .Y(n7069) );
  NAND2X1 U649 ( .A(arr[311]), .B(n2789), .Y(n4827) );
  OAI21X1 U650 ( .A(n4497), .B(n2788), .C(n4828), .Y(n7070) );
  NAND2X1 U651 ( .A(arr[312]), .B(n2789), .Y(n4828) );
  OAI21X1 U652 ( .A(n4499), .B(n2788), .C(n4829), .Y(n7071) );
  NAND2X1 U653 ( .A(arr[313]), .B(n2789), .Y(n4829) );
  OAI21X1 U654 ( .A(n4501), .B(n2787), .C(n4830), .Y(n7072) );
  NAND2X1 U655 ( .A(arr[314]), .B(n2789), .Y(n4830) );
  OAI21X1 U656 ( .A(n4503), .B(n2787), .C(n4831), .Y(n7073) );
  NAND2X1 U657 ( .A(arr[315]), .B(n2789), .Y(n4831) );
  OAI21X1 U658 ( .A(n4505), .B(n2787), .C(n4832), .Y(n7074) );
  NAND2X1 U659 ( .A(arr[316]), .B(n2789), .Y(n4832) );
  OAI21X1 U660 ( .A(n4507), .B(n2787), .C(n4833), .Y(n7075) );
  NAND2X1 U661 ( .A(arr[317]), .B(n2789), .Y(n4833) );
  OAI21X1 U662 ( .A(n4509), .B(n2787), .C(n4834), .Y(n7076) );
  NAND2X1 U663 ( .A(arr[318]), .B(n2789), .Y(n4834) );
  OAI21X1 U664 ( .A(n4511), .B(n2787), .C(n4835), .Y(n7077) );
  NAND2X1 U665 ( .A(arr[319]), .B(n2789), .Y(n4835) );
  OAI21X1 U666 ( .A(n4513), .B(n2789), .C(n4836), .Y(n7078) );
  NAND2X1 U667 ( .A(arr[320]), .B(n2789), .Y(n4836) );
  OAI21X1 U668 ( .A(n4515), .B(n2787), .C(n4837), .Y(n7079) );
  NAND2X1 U669 ( .A(arr[321]), .B(n2789), .Y(n4837) );
  OAI21X1 U670 ( .A(n4517), .B(n2788), .C(n4838), .Y(n7080) );
  NAND2X1 U671 ( .A(arr[322]), .B(n2789), .Y(n4838) );
  OAI21X1 U672 ( .A(n4519), .B(n2787), .C(n4839), .Y(n7081) );
  NAND2X1 U673 ( .A(arr[323]), .B(n2788), .Y(n4839) );
  OAI21X1 U674 ( .A(n4521), .B(n2788), .C(n4840), .Y(n7082) );
  NAND2X1 U675 ( .A(arr[324]), .B(n2789), .Y(n4840) );
  OAI21X1 U676 ( .A(n4523), .B(n2787), .C(n4841), .Y(n7083) );
  NAND2X1 U677 ( .A(arr[325]), .B(n2788), .Y(n4841) );
  OAI21X1 U678 ( .A(n4525), .B(n2787), .C(n4842), .Y(n7084) );
  NAND2X1 U679 ( .A(arr[326]), .B(n2789), .Y(n4842) );
  OAI21X1 U680 ( .A(n4527), .B(n2787), .C(n4843), .Y(n7085) );
  NAND2X1 U681 ( .A(arr[327]), .B(n2788), .Y(n4843) );
  OAI21X1 U682 ( .A(n4529), .B(n2787), .C(n4844), .Y(n7086) );
  NAND2X1 U683 ( .A(arr[328]), .B(n2788), .Y(n4844) );
  OAI21X1 U684 ( .A(n4531), .B(n2787), .C(n4845), .Y(n7087) );
  NAND2X1 U685 ( .A(arr[329]), .B(n2789), .Y(n4845) );
  OAI21X1 U687 ( .A(n4467), .B(n2784), .C(n4847), .Y(n7088) );
  NAND2X1 U688 ( .A(arr[330]), .B(n2786), .Y(n4847) );
  OAI21X1 U689 ( .A(n4469), .B(n2784), .C(n4848), .Y(n7089) );
  NAND2X1 U690 ( .A(arr[331]), .B(n2786), .Y(n4848) );
  OAI21X1 U691 ( .A(n4471), .B(n2784), .C(n4849), .Y(n7090) );
  NAND2X1 U692 ( .A(arr[332]), .B(n2786), .Y(n4849) );
  OAI21X1 U693 ( .A(n4473), .B(n2784), .C(n4850), .Y(n7091) );
  NAND2X1 U694 ( .A(arr[333]), .B(n2786), .Y(n4850) );
  OAI21X1 U695 ( .A(n4475), .B(n2785), .C(n4851), .Y(n7092) );
  NAND2X1 U696 ( .A(arr[334]), .B(n2786), .Y(n4851) );
  OAI21X1 U697 ( .A(n4477), .B(n2785), .C(n4852), .Y(n7093) );
  NAND2X1 U698 ( .A(arr[335]), .B(n2785), .Y(n4852) );
  OAI21X1 U699 ( .A(n4479), .B(n2785), .C(n4853), .Y(n7094) );
  NAND2X1 U700 ( .A(arr[336]), .B(n2786), .Y(n4853) );
  OAI21X1 U701 ( .A(n4481), .B(n2786), .C(n4854), .Y(n7095) );
  NAND2X1 U702 ( .A(arr[337]), .B(n2786), .Y(n4854) );
  OAI21X1 U703 ( .A(n4483), .B(n2785), .C(n4855), .Y(n7096) );
  NAND2X1 U704 ( .A(arr[338]), .B(n2786), .Y(n4855) );
  OAI21X1 U705 ( .A(n4485), .B(n2786), .C(n4856), .Y(n7097) );
  NAND2X1 U706 ( .A(arr[339]), .B(n2784), .Y(n4856) );
  OAI21X1 U707 ( .A(n4487), .B(n2786), .C(n4857), .Y(n7098) );
  NAND2X1 U708 ( .A(arr[340]), .B(n2786), .Y(n4857) );
  OAI21X1 U709 ( .A(n4489), .B(n2785), .C(n4858), .Y(n7099) );
  NAND2X1 U710 ( .A(arr[341]), .B(n2784), .Y(n4858) );
  OAI21X1 U711 ( .A(n4491), .B(n2786), .C(n4859), .Y(n7100) );
  NAND2X1 U712 ( .A(arr[342]), .B(n2785), .Y(n4859) );
  OAI21X1 U713 ( .A(n4493), .B(n2786), .C(n4860), .Y(n7101) );
  NAND2X1 U714 ( .A(arr[343]), .B(n2785), .Y(n4860) );
  OAI21X1 U715 ( .A(n4495), .B(n2785), .C(n4861), .Y(n7102) );
  NAND2X1 U716 ( .A(arr[344]), .B(n2786), .Y(n4861) );
  OAI21X1 U717 ( .A(n4497), .B(n2786), .C(n4862), .Y(n7103) );
  NAND2X1 U718 ( .A(arr[345]), .B(n2784), .Y(n4862) );
  OAI21X1 U719 ( .A(n4499), .B(n2786), .C(n4863), .Y(n7104) );
  NAND2X1 U720 ( .A(arr[346]), .B(n2786), .Y(n4863) );
  OAI21X1 U721 ( .A(n4501), .B(n2785), .C(n4864), .Y(n7105) );
  NAND2X1 U722 ( .A(arr[347]), .B(n2784), .Y(n4864) );
  OAI21X1 U723 ( .A(n4503), .B(n2785), .C(n4865), .Y(n7106) );
  NAND2X1 U724 ( .A(arr[348]), .B(n2785), .Y(n4865) );
  OAI21X1 U725 ( .A(n4505), .B(n2785), .C(n4866), .Y(n7107) );
  NAND2X1 U726 ( .A(arr[349]), .B(n2786), .Y(n4866) );
  OAI21X1 U727 ( .A(n4507), .B(n2785), .C(n4867), .Y(n7108) );
  NAND2X1 U728 ( .A(arr[350]), .B(n2784), .Y(n4867) );
  OAI21X1 U729 ( .A(n4509), .B(n2785), .C(n4868), .Y(n7109) );
  NAND2X1 U730 ( .A(arr[351]), .B(n2785), .Y(n4868) );
  OAI21X1 U731 ( .A(n4511), .B(n2785), .C(n4869), .Y(n7110) );
  NAND2X1 U732 ( .A(arr[352]), .B(n2786), .Y(n4869) );
  OAI21X1 U733 ( .A(n4513), .B(n2784), .C(n4870), .Y(n7111) );
  NAND2X1 U734 ( .A(arr[353]), .B(n2786), .Y(n4870) );
  OAI21X1 U735 ( .A(n4515), .B(n2785), .C(n4871), .Y(n7112) );
  NAND2X1 U736 ( .A(arr[354]), .B(n2786), .Y(n4871) );
  OAI21X1 U737 ( .A(n4517), .B(n2784), .C(n4872), .Y(n7113) );
  NAND2X1 U738 ( .A(arr[355]), .B(n2785), .Y(n4872) );
  OAI21X1 U739 ( .A(n4519), .B(n2784), .C(n4873), .Y(n7114) );
  NAND2X1 U740 ( .A(arr[356]), .B(n2784), .Y(n4873) );
  OAI21X1 U741 ( .A(n4521), .B(n2784), .C(n4874), .Y(n7115) );
  NAND2X1 U742 ( .A(arr[357]), .B(n2786), .Y(n4874) );
  OAI21X1 U743 ( .A(n4523), .B(n2784), .C(n4875), .Y(n7116) );
  NAND2X1 U744 ( .A(arr[358]), .B(n2785), .Y(n4875) );
  OAI21X1 U745 ( .A(n4525), .B(n2784), .C(n4876), .Y(n7117) );
  NAND2X1 U746 ( .A(arr[359]), .B(n2785), .Y(n4876) );
  OAI21X1 U747 ( .A(n4527), .B(n2784), .C(n4877), .Y(n7118) );
  NAND2X1 U748 ( .A(arr[360]), .B(n2784), .Y(n4877) );
  OAI21X1 U749 ( .A(n4529), .B(n2784), .C(n4878), .Y(n7119) );
  NAND2X1 U750 ( .A(arr[361]), .B(n2786), .Y(n4878) );
  OAI21X1 U751 ( .A(n4531), .B(n2784), .C(n4879), .Y(n7120) );
  NAND2X1 U752 ( .A(arr[362]), .B(n2784), .Y(n4879) );
  OAI21X1 U754 ( .A(n4467), .B(n2783), .C(n4882), .Y(n7121) );
  NAND2X1 U755 ( .A(arr[363]), .B(n2782), .Y(n4882) );
  OAI21X1 U756 ( .A(n4469), .B(n2781), .C(n4883), .Y(n7122) );
  NAND2X1 U757 ( .A(arr[364]), .B(n2782), .Y(n4883) );
  OAI21X1 U758 ( .A(n4471), .B(n2781), .C(n4884), .Y(n7123) );
  NAND2X1 U759 ( .A(arr[365]), .B(n2782), .Y(n4884) );
  OAI21X1 U760 ( .A(n4473), .B(n2781), .C(n4885), .Y(n7124) );
  NAND2X1 U761 ( .A(arr[366]), .B(n2782), .Y(n4885) );
  OAI21X1 U762 ( .A(n4475), .B(n2781), .C(n4886), .Y(n7125) );
  NAND2X1 U763 ( .A(arr[367]), .B(n2782), .Y(n4886) );
  OAI21X1 U764 ( .A(n4477), .B(n2781), .C(n4887), .Y(n7126) );
  NAND2X1 U765 ( .A(arr[368]), .B(n2783), .Y(n4887) );
  OAI21X1 U766 ( .A(n4479), .B(n2781), .C(n4888), .Y(n7127) );
  NAND2X1 U767 ( .A(arr[369]), .B(n2783), .Y(n4888) );
  OAI21X1 U768 ( .A(n4481), .B(n2782), .C(n4889), .Y(n7128) );
  NAND2X1 U769 ( .A(arr[370]), .B(n2782), .Y(n4889) );
  OAI21X1 U770 ( .A(n4483), .B(n2781), .C(n4890), .Y(n7129) );
  NAND2X1 U771 ( .A(arr[371]), .B(n2782), .Y(n4890) );
  OAI21X1 U772 ( .A(n4485), .B(n2782), .C(n4891), .Y(n7130) );
  NAND2X1 U773 ( .A(arr[372]), .B(n2783), .Y(n4891) );
  OAI21X1 U774 ( .A(n4487), .B(n2782), .C(n4892), .Y(n7131) );
  NAND2X1 U775 ( .A(arr[373]), .B(n2783), .Y(n4892) );
  OAI21X1 U776 ( .A(n4489), .B(n2781), .C(n4893), .Y(n7132) );
  NAND2X1 U777 ( .A(arr[374]), .B(n2783), .Y(n4893) );
  OAI21X1 U778 ( .A(n4491), .B(n2782), .C(n4894), .Y(n7133) );
  NAND2X1 U779 ( .A(arr[375]), .B(n2783), .Y(n4894) );
  OAI21X1 U780 ( .A(n4493), .B(n2782), .C(n4895), .Y(n7134) );
  NAND2X1 U781 ( .A(arr[376]), .B(n2783), .Y(n4895) );
  OAI21X1 U782 ( .A(n4495), .B(n2781), .C(n4896), .Y(n7135) );
  NAND2X1 U783 ( .A(arr[377]), .B(n2783), .Y(n4896) );
  OAI21X1 U784 ( .A(n4497), .B(n2782), .C(n4897), .Y(n7136) );
  NAND2X1 U785 ( .A(arr[378]), .B(n2783), .Y(n4897) );
  OAI21X1 U786 ( .A(n4499), .B(n2782), .C(n4898), .Y(n7137) );
  NAND2X1 U787 ( .A(arr[379]), .B(n2783), .Y(n4898) );
  OAI21X1 U788 ( .A(n4501), .B(n2781), .C(n4899), .Y(n7138) );
  NAND2X1 U789 ( .A(arr[380]), .B(n2783), .Y(n4899) );
  OAI21X1 U790 ( .A(n4503), .B(n2781), .C(n4900), .Y(n7139) );
  NAND2X1 U791 ( .A(arr[381]), .B(n2783), .Y(n4900) );
  OAI21X1 U792 ( .A(n4505), .B(n2781), .C(n4901), .Y(n7140) );
  NAND2X1 U793 ( .A(arr[382]), .B(n2783), .Y(n4901) );
  OAI21X1 U794 ( .A(n4507), .B(n2781), .C(n4902), .Y(n7141) );
  NAND2X1 U795 ( .A(arr[383]), .B(n2783), .Y(n4902) );
  OAI21X1 U796 ( .A(n4509), .B(n2781), .C(n4903), .Y(n7142) );
  NAND2X1 U797 ( .A(arr[384]), .B(n2783), .Y(n4903) );
  OAI21X1 U798 ( .A(n4511), .B(n2781), .C(n4904), .Y(n7143) );
  NAND2X1 U799 ( .A(arr[385]), .B(n2783), .Y(n4904) );
  OAI21X1 U800 ( .A(n4513), .B(n2783), .C(n4905), .Y(n7144) );
  NAND2X1 U801 ( .A(arr[386]), .B(n2783), .Y(n4905) );
  OAI21X1 U802 ( .A(n4515), .B(n2781), .C(n4906), .Y(n7145) );
  NAND2X1 U803 ( .A(arr[387]), .B(n2783), .Y(n4906) );
  OAI21X1 U804 ( .A(n4517), .B(n2782), .C(n4907), .Y(n7146) );
  NAND2X1 U805 ( .A(arr[388]), .B(n2783), .Y(n4907) );
  OAI21X1 U806 ( .A(n4519), .B(n2781), .C(n4908), .Y(n7147) );
  NAND2X1 U807 ( .A(arr[389]), .B(n2782), .Y(n4908) );
  OAI21X1 U808 ( .A(n4521), .B(n2782), .C(n4909), .Y(n7148) );
  NAND2X1 U809 ( .A(arr[390]), .B(n2783), .Y(n4909) );
  OAI21X1 U810 ( .A(n4523), .B(n2781), .C(n4910), .Y(n7149) );
  NAND2X1 U811 ( .A(arr[391]), .B(n2782), .Y(n4910) );
  OAI21X1 U812 ( .A(n4525), .B(n2781), .C(n4911), .Y(n7150) );
  NAND2X1 U813 ( .A(arr[392]), .B(n2783), .Y(n4911) );
  OAI21X1 U814 ( .A(n4527), .B(n2781), .C(n4912), .Y(n7151) );
  NAND2X1 U815 ( .A(arr[393]), .B(n2782), .Y(n4912) );
  OAI21X1 U816 ( .A(n4529), .B(n2781), .C(n4913), .Y(n7152) );
  NAND2X1 U817 ( .A(arr[394]), .B(n2782), .Y(n4913) );
  OAI21X1 U818 ( .A(n4531), .B(n2781), .C(n4914), .Y(n7153) );
  NAND2X1 U819 ( .A(arr[395]), .B(n2783), .Y(n4914) );
  OAI21X1 U821 ( .A(n4467), .B(n2778), .C(n4916), .Y(n7154) );
  NAND2X1 U822 ( .A(arr[396]), .B(n2780), .Y(n4916) );
  OAI21X1 U823 ( .A(n4469), .B(n2778), .C(n4917), .Y(n7155) );
  NAND2X1 U824 ( .A(arr[397]), .B(n2780), .Y(n4917) );
  OAI21X1 U825 ( .A(n4471), .B(n2778), .C(n4918), .Y(n7156) );
  NAND2X1 U826 ( .A(arr[398]), .B(n2780), .Y(n4918) );
  OAI21X1 U827 ( .A(n4473), .B(n2778), .C(n4919), .Y(n7157) );
  NAND2X1 U828 ( .A(arr[399]), .B(n2780), .Y(n4919) );
  OAI21X1 U829 ( .A(n4475), .B(n2779), .C(n4920), .Y(n7158) );
  NAND2X1 U830 ( .A(arr[400]), .B(n2780), .Y(n4920) );
  OAI21X1 U831 ( .A(n4477), .B(n2779), .C(n4921), .Y(n7159) );
  NAND2X1 U832 ( .A(arr[401]), .B(n2779), .Y(n4921) );
  OAI21X1 U833 ( .A(n4479), .B(n2779), .C(n4922), .Y(n7160) );
  NAND2X1 U834 ( .A(arr[402]), .B(n2780), .Y(n4922) );
  OAI21X1 U835 ( .A(n4481), .B(n2780), .C(n4923), .Y(n7161) );
  NAND2X1 U836 ( .A(arr[403]), .B(n2780), .Y(n4923) );
  OAI21X1 U837 ( .A(n4483), .B(n2779), .C(n4924), .Y(n7162) );
  NAND2X1 U838 ( .A(arr[404]), .B(n2780), .Y(n4924) );
  OAI21X1 U839 ( .A(n4485), .B(n2780), .C(n4925), .Y(n7163) );
  NAND2X1 U840 ( .A(arr[405]), .B(n2778), .Y(n4925) );
  OAI21X1 U841 ( .A(n4487), .B(n2780), .C(n4926), .Y(n7164) );
  NAND2X1 U842 ( .A(arr[406]), .B(n2780), .Y(n4926) );
  OAI21X1 U843 ( .A(n4489), .B(n2779), .C(n4927), .Y(n7165) );
  NAND2X1 U844 ( .A(arr[407]), .B(n2778), .Y(n4927) );
  OAI21X1 U845 ( .A(n4491), .B(n2780), .C(n4928), .Y(n7166) );
  NAND2X1 U846 ( .A(arr[408]), .B(n2779), .Y(n4928) );
  OAI21X1 U847 ( .A(n4493), .B(n2780), .C(n4929), .Y(n7167) );
  NAND2X1 U848 ( .A(arr[409]), .B(n2779), .Y(n4929) );
  OAI21X1 U849 ( .A(n4495), .B(n2779), .C(n4930), .Y(n7168) );
  NAND2X1 U850 ( .A(arr[410]), .B(n2780), .Y(n4930) );
  OAI21X1 U851 ( .A(n4497), .B(n2780), .C(n4931), .Y(n7169) );
  NAND2X1 U852 ( .A(arr[411]), .B(n2778), .Y(n4931) );
  OAI21X1 U853 ( .A(n4499), .B(n2780), .C(n4932), .Y(n7170) );
  NAND2X1 U854 ( .A(arr[412]), .B(n2780), .Y(n4932) );
  OAI21X1 U855 ( .A(n4501), .B(n2779), .C(n4933), .Y(n7171) );
  NAND2X1 U856 ( .A(arr[413]), .B(n2778), .Y(n4933) );
  OAI21X1 U857 ( .A(n4503), .B(n2779), .C(n4934), .Y(n7172) );
  NAND2X1 U858 ( .A(arr[414]), .B(n2779), .Y(n4934) );
  OAI21X1 U859 ( .A(n4505), .B(n2779), .C(n4935), .Y(n7173) );
  NAND2X1 U860 ( .A(arr[415]), .B(n2780), .Y(n4935) );
  OAI21X1 U861 ( .A(n4507), .B(n2779), .C(n4936), .Y(n7174) );
  NAND2X1 U862 ( .A(arr[416]), .B(n2778), .Y(n4936) );
  OAI21X1 U863 ( .A(n4509), .B(n2779), .C(n4937), .Y(n7175) );
  NAND2X1 U864 ( .A(arr[417]), .B(n2779), .Y(n4937) );
  OAI21X1 U865 ( .A(n4511), .B(n2779), .C(n4938), .Y(n7176) );
  NAND2X1 U866 ( .A(arr[418]), .B(n2780), .Y(n4938) );
  OAI21X1 U867 ( .A(n4513), .B(n2778), .C(n4939), .Y(n7177) );
  NAND2X1 U868 ( .A(arr[419]), .B(n2780), .Y(n4939) );
  OAI21X1 U869 ( .A(n4515), .B(n2779), .C(n4940), .Y(n7178) );
  NAND2X1 U870 ( .A(arr[420]), .B(n2780), .Y(n4940) );
  OAI21X1 U871 ( .A(n4517), .B(n2778), .C(n4941), .Y(n7179) );
  NAND2X1 U872 ( .A(arr[421]), .B(n2779), .Y(n4941) );
  OAI21X1 U873 ( .A(n4519), .B(n2778), .C(n4942), .Y(n7180) );
  NAND2X1 U874 ( .A(arr[422]), .B(n2778), .Y(n4942) );
  OAI21X1 U875 ( .A(n4521), .B(n2778), .C(n4943), .Y(n7181) );
  NAND2X1 U876 ( .A(arr[423]), .B(n2780), .Y(n4943) );
  OAI21X1 U877 ( .A(n4523), .B(n2778), .C(n4944), .Y(n7182) );
  NAND2X1 U878 ( .A(arr[424]), .B(n2779), .Y(n4944) );
  OAI21X1 U879 ( .A(n4525), .B(n2778), .C(n4945), .Y(n7183) );
  NAND2X1 U880 ( .A(arr[425]), .B(n2779), .Y(n4945) );
  OAI21X1 U881 ( .A(n4527), .B(n2778), .C(n4946), .Y(n7184) );
  NAND2X1 U882 ( .A(arr[426]), .B(n2778), .Y(n4946) );
  OAI21X1 U883 ( .A(n4529), .B(n2778), .C(n4947), .Y(n7185) );
  NAND2X1 U884 ( .A(arr[427]), .B(n2780), .Y(n4947) );
  OAI21X1 U885 ( .A(n4531), .B(n2778), .C(n4948), .Y(n7186) );
  NAND2X1 U886 ( .A(arr[428]), .B(n2778), .Y(n4948) );
  OAI21X1 U888 ( .A(n4467), .B(n2777), .C(n4951), .Y(n7187) );
  NAND2X1 U889 ( .A(arr[429]), .B(n2776), .Y(n4951) );
  OAI21X1 U890 ( .A(n4469), .B(n2775), .C(n4952), .Y(n7188) );
  NAND2X1 U891 ( .A(arr[430]), .B(n2776), .Y(n4952) );
  OAI21X1 U892 ( .A(n4471), .B(n2775), .C(n4953), .Y(n7189) );
  NAND2X1 U893 ( .A(arr[431]), .B(n2776), .Y(n4953) );
  OAI21X1 U894 ( .A(n4473), .B(n2775), .C(n4954), .Y(n7190) );
  NAND2X1 U895 ( .A(arr[432]), .B(n2776), .Y(n4954) );
  OAI21X1 U896 ( .A(n4475), .B(n2775), .C(n4955), .Y(n7191) );
  NAND2X1 U897 ( .A(arr[433]), .B(n2776), .Y(n4955) );
  OAI21X1 U898 ( .A(n4477), .B(n2775), .C(n4956), .Y(n7192) );
  NAND2X1 U899 ( .A(arr[434]), .B(n2777), .Y(n4956) );
  OAI21X1 U900 ( .A(n4479), .B(n2775), .C(n4957), .Y(n7193) );
  NAND2X1 U901 ( .A(arr[435]), .B(n2777), .Y(n4957) );
  OAI21X1 U902 ( .A(n4481), .B(n2776), .C(n4958), .Y(n7194) );
  NAND2X1 U903 ( .A(arr[436]), .B(n2776), .Y(n4958) );
  OAI21X1 U904 ( .A(n4483), .B(n2775), .C(n4959), .Y(n7195) );
  NAND2X1 U905 ( .A(arr[437]), .B(n2776), .Y(n4959) );
  OAI21X1 U906 ( .A(n4485), .B(n2776), .C(n4960), .Y(n7196) );
  NAND2X1 U907 ( .A(arr[438]), .B(n2777), .Y(n4960) );
  OAI21X1 U908 ( .A(n4487), .B(n2776), .C(n4961), .Y(n7197) );
  NAND2X1 U909 ( .A(arr[439]), .B(n2777), .Y(n4961) );
  OAI21X1 U910 ( .A(n4489), .B(n2775), .C(n4962), .Y(n7198) );
  NAND2X1 U911 ( .A(arr[440]), .B(n2777), .Y(n4962) );
  OAI21X1 U912 ( .A(n4491), .B(n2776), .C(n4963), .Y(n7199) );
  NAND2X1 U913 ( .A(arr[441]), .B(n2777), .Y(n4963) );
  OAI21X1 U914 ( .A(n4493), .B(n2776), .C(n4964), .Y(n7200) );
  NAND2X1 U915 ( .A(arr[442]), .B(n2777), .Y(n4964) );
  OAI21X1 U916 ( .A(n4495), .B(n2775), .C(n4965), .Y(n7201) );
  NAND2X1 U917 ( .A(arr[443]), .B(n2777), .Y(n4965) );
  OAI21X1 U918 ( .A(n4497), .B(n2776), .C(n4966), .Y(n7202) );
  NAND2X1 U919 ( .A(arr[444]), .B(n2777), .Y(n4966) );
  OAI21X1 U920 ( .A(n4499), .B(n2776), .C(n4967), .Y(n7203) );
  NAND2X1 U921 ( .A(arr[445]), .B(n2777), .Y(n4967) );
  OAI21X1 U922 ( .A(n4501), .B(n2775), .C(n4968), .Y(n7204) );
  NAND2X1 U923 ( .A(arr[446]), .B(n2777), .Y(n4968) );
  OAI21X1 U924 ( .A(n4503), .B(n2775), .C(n4969), .Y(n7205) );
  NAND2X1 U925 ( .A(arr[447]), .B(n2777), .Y(n4969) );
  OAI21X1 U926 ( .A(n4505), .B(n2775), .C(n4970), .Y(n7206) );
  NAND2X1 U927 ( .A(arr[448]), .B(n2777), .Y(n4970) );
  OAI21X1 U928 ( .A(n4507), .B(n2775), .C(n4971), .Y(n7207) );
  NAND2X1 U929 ( .A(arr[449]), .B(n2777), .Y(n4971) );
  OAI21X1 U930 ( .A(n4509), .B(n2775), .C(n4972), .Y(n7208) );
  NAND2X1 U931 ( .A(arr[450]), .B(n2777), .Y(n4972) );
  OAI21X1 U932 ( .A(n4511), .B(n2775), .C(n4973), .Y(n7209) );
  NAND2X1 U933 ( .A(arr[451]), .B(n2777), .Y(n4973) );
  OAI21X1 U934 ( .A(n4513), .B(n2777), .C(n4974), .Y(n7210) );
  NAND2X1 U935 ( .A(arr[452]), .B(n2777), .Y(n4974) );
  OAI21X1 U936 ( .A(n4515), .B(n2775), .C(n4975), .Y(n7211) );
  NAND2X1 U937 ( .A(arr[453]), .B(n2777), .Y(n4975) );
  OAI21X1 U938 ( .A(n4517), .B(n2776), .C(n4976), .Y(n7212) );
  NAND2X1 U939 ( .A(arr[454]), .B(n2777), .Y(n4976) );
  OAI21X1 U940 ( .A(n4519), .B(n2775), .C(n4977), .Y(n7213) );
  NAND2X1 U941 ( .A(arr[455]), .B(n2776), .Y(n4977) );
  OAI21X1 U942 ( .A(n4521), .B(n2776), .C(n4978), .Y(n7214) );
  NAND2X1 U943 ( .A(arr[456]), .B(n2777), .Y(n4978) );
  OAI21X1 U944 ( .A(n4523), .B(n2775), .C(n4979), .Y(n7215) );
  NAND2X1 U945 ( .A(arr[457]), .B(n2776), .Y(n4979) );
  OAI21X1 U946 ( .A(n4525), .B(n2775), .C(n4980), .Y(n7216) );
  NAND2X1 U947 ( .A(arr[458]), .B(n2777), .Y(n4980) );
  OAI21X1 U948 ( .A(n4527), .B(n2775), .C(n4981), .Y(n7217) );
  NAND2X1 U949 ( .A(arr[459]), .B(n2776), .Y(n4981) );
  OAI21X1 U950 ( .A(n4529), .B(n2775), .C(n4982), .Y(n7218) );
  NAND2X1 U951 ( .A(arr[460]), .B(n2776), .Y(n4982) );
  OAI21X1 U952 ( .A(n4531), .B(n2775), .C(n4983), .Y(n7219) );
  NAND2X1 U953 ( .A(arr[461]), .B(n2777), .Y(n4983) );
  OAI21X1 U955 ( .A(n4467), .B(n2772), .C(n4985), .Y(n7220) );
  NAND2X1 U956 ( .A(arr[462]), .B(n2774), .Y(n4985) );
  OAI21X1 U957 ( .A(n4469), .B(n2772), .C(n4986), .Y(n7221) );
  NAND2X1 U958 ( .A(arr[463]), .B(n2774), .Y(n4986) );
  OAI21X1 U959 ( .A(n4471), .B(n2772), .C(n4987), .Y(n7222) );
  NAND2X1 U960 ( .A(arr[464]), .B(n2774), .Y(n4987) );
  OAI21X1 U961 ( .A(n4473), .B(n2772), .C(n4988), .Y(n7223) );
  NAND2X1 U962 ( .A(arr[465]), .B(n2774), .Y(n4988) );
  OAI21X1 U963 ( .A(n4475), .B(n2773), .C(n4989), .Y(n7224) );
  NAND2X1 U964 ( .A(arr[466]), .B(n2774), .Y(n4989) );
  OAI21X1 U965 ( .A(n4477), .B(n2773), .C(n4990), .Y(n7225) );
  NAND2X1 U966 ( .A(arr[467]), .B(n2773), .Y(n4990) );
  OAI21X1 U967 ( .A(n4479), .B(n2773), .C(n4991), .Y(n7226) );
  NAND2X1 U968 ( .A(arr[468]), .B(n2774), .Y(n4991) );
  OAI21X1 U969 ( .A(n4481), .B(n2774), .C(n4992), .Y(n7227) );
  NAND2X1 U970 ( .A(arr[469]), .B(n2774), .Y(n4992) );
  OAI21X1 U971 ( .A(n4483), .B(n2773), .C(n4993), .Y(n7228) );
  NAND2X1 U972 ( .A(arr[470]), .B(n2774), .Y(n4993) );
  OAI21X1 U973 ( .A(n4485), .B(n2774), .C(n4994), .Y(n7229) );
  NAND2X1 U974 ( .A(arr[471]), .B(n2772), .Y(n4994) );
  OAI21X1 U975 ( .A(n4487), .B(n2774), .C(n4995), .Y(n7230) );
  NAND2X1 U976 ( .A(arr[472]), .B(n2774), .Y(n4995) );
  OAI21X1 U977 ( .A(n4489), .B(n2773), .C(n4996), .Y(n7231) );
  NAND2X1 U978 ( .A(arr[473]), .B(n2772), .Y(n4996) );
  OAI21X1 U979 ( .A(n4491), .B(n2774), .C(n4997), .Y(n7232) );
  NAND2X1 U980 ( .A(arr[474]), .B(n2773), .Y(n4997) );
  OAI21X1 U981 ( .A(n4493), .B(n2774), .C(n4998), .Y(n7233) );
  NAND2X1 U982 ( .A(arr[475]), .B(n2773), .Y(n4998) );
  OAI21X1 U983 ( .A(n4495), .B(n2773), .C(n4999), .Y(n7234) );
  NAND2X1 U984 ( .A(arr[476]), .B(n2774), .Y(n4999) );
  OAI21X1 U985 ( .A(n4497), .B(n2774), .C(n5000), .Y(n7235) );
  NAND2X1 U986 ( .A(arr[477]), .B(n2772), .Y(n5000) );
  OAI21X1 U987 ( .A(n4499), .B(n2774), .C(n5001), .Y(n7236) );
  NAND2X1 U988 ( .A(arr[478]), .B(n2774), .Y(n5001) );
  OAI21X1 U989 ( .A(n4501), .B(n2773), .C(n5002), .Y(n7237) );
  NAND2X1 U990 ( .A(arr[479]), .B(n2772), .Y(n5002) );
  OAI21X1 U991 ( .A(n4503), .B(n2773), .C(n5003), .Y(n7238) );
  NAND2X1 U992 ( .A(arr[480]), .B(n2773), .Y(n5003) );
  OAI21X1 U993 ( .A(n4505), .B(n2773), .C(n5004), .Y(n7239) );
  NAND2X1 U994 ( .A(arr[481]), .B(n2774), .Y(n5004) );
  OAI21X1 U995 ( .A(n4507), .B(n2773), .C(n5005), .Y(n7240) );
  NAND2X1 U996 ( .A(arr[482]), .B(n2772), .Y(n5005) );
  OAI21X1 U997 ( .A(n4509), .B(n2773), .C(n5006), .Y(n7241) );
  NAND2X1 U998 ( .A(arr[483]), .B(n2773), .Y(n5006) );
  OAI21X1 U999 ( .A(n4511), .B(n2773), .C(n5007), .Y(n7242) );
  NAND2X1 U1000 ( .A(arr[484]), .B(n2774), .Y(n5007) );
  OAI21X1 U1001 ( .A(n4513), .B(n2772), .C(n5008), .Y(n7243) );
  NAND2X1 U1002 ( .A(arr[485]), .B(n2774), .Y(n5008) );
  OAI21X1 U1003 ( .A(n4515), .B(n2773), .C(n5009), .Y(n7244) );
  NAND2X1 U1004 ( .A(arr[486]), .B(n2774), .Y(n5009) );
  OAI21X1 U1005 ( .A(n4517), .B(n2772), .C(n5010), .Y(n7245) );
  NAND2X1 U1006 ( .A(arr[487]), .B(n2773), .Y(n5010) );
  OAI21X1 U1007 ( .A(n4519), .B(n2772), .C(n5011), .Y(n7246) );
  NAND2X1 U1008 ( .A(arr[488]), .B(n2772), .Y(n5011) );
  OAI21X1 U1009 ( .A(n4521), .B(n2772), .C(n5012), .Y(n7247) );
  NAND2X1 U1010 ( .A(arr[489]), .B(n2774), .Y(n5012) );
  OAI21X1 U1011 ( .A(n4523), .B(n2772), .C(n5013), .Y(n7248) );
  NAND2X1 U1012 ( .A(arr[490]), .B(n2773), .Y(n5013) );
  OAI21X1 U1013 ( .A(n4525), .B(n2772), .C(n5014), .Y(n7249) );
  NAND2X1 U1014 ( .A(arr[491]), .B(n2773), .Y(n5014) );
  OAI21X1 U1015 ( .A(n4527), .B(n2772), .C(n5015), .Y(n7250) );
  NAND2X1 U1016 ( .A(arr[492]), .B(n2772), .Y(n5015) );
  OAI21X1 U1017 ( .A(n4529), .B(n2772), .C(n5016), .Y(n7251) );
  NAND2X1 U1018 ( .A(arr[493]), .B(n2774), .Y(n5016) );
  OAI21X1 U1019 ( .A(n4531), .B(n2772), .C(n5017), .Y(n7252) );
  NAND2X1 U1020 ( .A(arr[494]), .B(n2772), .Y(n5017) );
  OAI21X1 U1022 ( .A(n4467), .B(n2771), .C(n5020), .Y(n7253) );
  NAND2X1 U1023 ( .A(arr[495]), .B(n2770), .Y(n5020) );
  OAI21X1 U1024 ( .A(n4469), .B(n2769), .C(n5021), .Y(n7254) );
  NAND2X1 U1025 ( .A(arr[496]), .B(n2770), .Y(n5021) );
  OAI21X1 U1026 ( .A(n4471), .B(n2769), .C(n5022), .Y(n7255) );
  NAND2X1 U1027 ( .A(arr[497]), .B(n2770), .Y(n5022) );
  OAI21X1 U1028 ( .A(n4473), .B(n2769), .C(n5023), .Y(n7256) );
  NAND2X1 U1029 ( .A(arr[498]), .B(n2770), .Y(n5023) );
  OAI21X1 U1030 ( .A(n4475), .B(n2769), .C(n5024), .Y(n7257) );
  NAND2X1 U1031 ( .A(arr[499]), .B(n2770), .Y(n5024) );
  OAI21X1 U1032 ( .A(n4477), .B(n2769), .C(n5025), .Y(n7258) );
  NAND2X1 U1033 ( .A(arr[500]), .B(n2771), .Y(n5025) );
  OAI21X1 U1034 ( .A(n4479), .B(n2769), .C(n5026), .Y(n7259) );
  NAND2X1 U1035 ( .A(arr[501]), .B(n2771), .Y(n5026) );
  OAI21X1 U1036 ( .A(n4481), .B(n2770), .C(n5027), .Y(n7260) );
  NAND2X1 U1037 ( .A(arr[502]), .B(n2770), .Y(n5027) );
  OAI21X1 U1038 ( .A(n4483), .B(n2769), .C(n5028), .Y(n7261) );
  NAND2X1 U1039 ( .A(arr[503]), .B(n2770), .Y(n5028) );
  OAI21X1 U1040 ( .A(n4485), .B(n2770), .C(n5029), .Y(n7262) );
  NAND2X1 U1041 ( .A(arr[504]), .B(n2771), .Y(n5029) );
  OAI21X1 U1042 ( .A(n4487), .B(n2770), .C(n5030), .Y(n7263) );
  NAND2X1 U1043 ( .A(arr[505]), .B(n2771), .Y(n5030) );
  OAI21X1 U1044 ( .A(n4489), .B(n2769), .C(n5031), .Y(n7264) );
  NAND2X1 U1045 ( .A(arr[506]), .B(n2771), .Y(n5031) );
  OAI21X1 U1046 ( .A(n4491), .B(n2770), .C(n5032), .Y(n7265) );
  NAND2X1 U1047 ( .A(arr[507]), .B(n2771), .Y(n5032) );
  OAI21X1 U1048 ( .A(n4493), .B(n2770), .C(n5033), .Y(n7266) );
  NAND2X1 U1049 ( .A(arr[508]), .B(n2771), .Y(n5033) );
  OAI21X1 U1050 ( .A(n4495), .B(n2769), .C(n5034), .Y(n7267) );
  NAND2X1 U1051 ( .A(arr[509]), .B(n2771), .Y(n5034) );
  OAI21X1 U1052 ( .A(n4497), .B(n2770), .C(n5035), .Y(n7268) );
  NAND2X1 U1053 ( .A(arr[510]), .B(n2771), .Y(n5035) );
  OAI21X1 U1054 ( .A(n4499), .B(n2770), .C(n5036), .Y(n7269) );
  NAND2X1 U1055 ( .A(arr[511]), .B(n2771), .Y(n5036) );
  OAI21X1 U1056 ( .A(n4501), .B(n2769), .C(n5037), .Y(n7270) );
  NAND2X1 U1057 ( .A(arr[512]), .B(n2771), .Y(n5037) );
  OAI21X1 U1058 ( .A(n4503), .B(n2769), .C(n5038), .Y(n7271) );
  NAND2X1 U1059 ( .A(arr[513]), .B(n2771), .Y(n5038) );
  OAI21X1 U1060 ( .A(n4505), .B(n2769), .C(n5039), .Y(n7272) );
  NAND2X1 U1061 ( .A(arr[514]), .B(n2771), .Y(n5039) );
  OAI21X1 U1062 ( .A(n4507), .B(n2769), .C(n5040), .Y(n7273) );
  NAND2X1 U1063 ( .A(arr[515]), .B(n2771), .Y(n5040) );
  OAI21X1 U1064 ( .A(n4509), .B(n2769), .C(n5041), .Y(n7274) );
  NAND2X1 U1065 ( .A(arr[516]), .B(n2771), .Y(n5041) );
  OAI21X1 U1066 ( .A(n4511), .B(n2769), .C(n5042), .Y(n7275) );
  NAND2X1 U1067 ( .A(arr[517]), .B(n2771), .Y(n5042) );
  OAI21X1 U1068 ( .A(n4513), .B(n2771), .C(n5043), .Y(n7276) );
  NAND2X1 U1069 ( .A(arr[518]), .B(n2771), .Y(n5043) );
  OAI21X1 U1070 ( .A(n4515), .B(n2769), .C(n5044), .Y(n7277) );
  NAND2X1 U1071 ( .A(arr[519]), .B(n2771), .Y(n5044) );
  OAI21X1 U1072 ( .A(n4517), .B(n2770), .C(n5045), .Y(n7278) );
  NAND2X1 U1073 ( .A(arr[520]), .B(n2771), .Y(n5045) );
  OAI21X1 U1074 ( .A(n4519), .B(n2769), .C(n5046), .Y(n7279) );
  NAND2X1 U1075 ( .A(arr[521]), .B(n2770), .Y(n5046) );
  OAI21X1 U1076 ( .A(n4521), .B(n2770), .C(n5047), .Y(n7280) );
  NAND2X1 U1077 ( .A(arr[522]), .B(n2771), .Y(n5047) );
  OAI21X1 U1078 ( .A(n4523), .B(n2769), .C(n5048), .Y(n7281) );
  NAND2X1 U1079 ( .A(arr[523]), .B(n2770), .Y(n5048) );
  OAI21X1 U1080 ( .A(n4525), .B(n2769), .C(n5049), .Y(n7282) );
  NAND2X1 U1081 ( .A(arr[524]), .B(n2771), .Y(n5049) );
  OAI21X1 U1082 ( .A(n4527), .B(n2769), .C(n5050), .Y(n7283) );
  NAND2X1 U1083 ( .A(arr[525]), .B(n2770), .Y(n5050) );
  OAI21X1 U1084 ( .A(n4529), .B(n2769), .C(n5051), .Y(n7284) );
  NAND2X1 U1085 ( .A(arr[526]), .B(n2770), .Y(n5051) );
  OAI21X1 U1086 ( .A(n4531), .B(n2769), .C(n5052), .Y(n7285) );
  NAND2X1 U1087 ( .A(arr[527]), .B(n2771), .Y(n5052) );
  OAI21X1 U1089 ( .A(n4467), .B(n2766), .C(n5054), .Y(n7286) );
  NAND2X1 U1090 ( .A(arr[528]), .B(n2768), .Y(n5054) );
  OAI21X1 U1091 ( .A(n4469), .B(n2766), .C(n5055), .Y(n7287) );
  NAND2X1 U1092 ( .A(arr[529]), .B(n2768), .Y(n5055) );
  OAI21X1 U1093 ( .A(n4471), .B(n2766), .C(n5056), .Y(n7288) );
  NAND2X1 U1094 ( .A(arr[530]), .B(n2768), .Y(n5056) );
  OAI21X1 U1095 ( .A(n4473), .B(n2766), .C(n5057), .Y(n7289) );
  NAND2X1 U1096 ( .A(arr[531]), .B(n2768), .Y(n5057) );
  OAI21X1 U1097 ( .A(n4475), .B(n2767), .C(n5058), .Y(n7290) );
  NAND2X1 U1098 ( .A(arr[532]), .B(n2768), .Y(n5058) );
  OAI21X1 U1099 ( .A(n4477), .B(n2767), .C(n5059), .Y(n7291) );
  NAND2X1 U1100 ( .A(arr[533]), .B(n2767), .Y(n5059) );
  OAI21X1 U1101 ( .A(n4479), .B(n2767), .C(n5060), .Y(n7292) );
  NAND2X1 U1102 ( .A(arr[534]), .B(n2768), .Y(n5060) );
  OAI21X1 U1103 ( .A(n4481), .B(n2768), .C(n5061), .Y(n7293) );
  NAND2X1 U1104 ( .A(arr[535]), .B(n2768), .Y(n5061) );
  OAI21X1 U1105 ( .A(n4483), .B(n2767), .C(n5062), .Y(n7294) );
  NAND2X1 U1106 ( .A(arr[536]), .B(n2768), .Y(n5062) );
  OAI21X1 U1107 ( .A(n4485), .B(n2768), .C(n5063), .Y(n7295) );
  NAND2X1 U1108 ( .A(arr[537]), .B(n2766), .Y(n5063) );
  OAI21X1 U1109 ( .A(n4487), .B(n2768), .C(n5064), .Y(n7296) );
  NAND2X1 U1110 ( .A(arr[538]), .B(n2768), .Y(n5064) );
  OAI21X1 U1111 ( .A(n4489), .B(n2767), .C(n5065), .Y(n7297) );
  NAND2X1 U1112 ( .A(arr[539]), .B(n2766), .Y(n5065) );
  OAI21X1 U1113 ( .A(n4491), .B(n2768), .C(n5066), .Y(n7298) );
  NAND2X1 U1114 ( .A(arr[540]), .B(n2767), .Y(n5066) );
  OAI21X1 U1115 ( .A(n4493), .B(n2768), .C(n5067), .Y(n7299) );
  NAND2X1 U1116 ( .A(arr[541]), .B(n2767), .Y(n5067) );
  OAI21X1 U1117 ( .A(n4495), .B(n2767), .C(n5068), .Y(n7300) );
  NAND2X1 U1118 ( .A(arr[542]), .B(n2768), .Y(n5068) );
  OAI21X1 U1119 ( .A(n4497), .B(n2768), .C(n5069), .Y(n7301) );
  NAND2X1 U1120 ( .A(arr[543]), .B(n2766), .Y(n5069) );
  OAI21X1 U1121 ( .A(n4499), .B(n2768), .C(n5070), .Y(n7302) );
  NAND2X1 U1122 ( .A(arr[544]), .B(n2768), .Y(n5070) );
  OAI21X1 U1123 ( .A(n4501), .B(n2767), .C(n5071), .Y(n7303) );
  NAND2X1 U1124 ( .A(arr[545]), .B(n2766), .Y(n5071) );
  OAI21X1 U1125 ( .A(n4503), .B(n2767), .C(n5072), .Y(n7304) );
  NAND2X1 U1126 ( .A(arr[546]), .B(n2767), .Y(n5072) );
  OAI21X1 U1127 ( .A(n4505), .B(n2767), .C(n5073), .Y(n7305) );
  NAND2X1 U1128 ( .A(arr[547]), .B(n2768), .Y(n5073) );
  OAI21X1 U1129 ( .A(n4507), .B(n2767), .C(n5074), .Y(n7306) );
  NAND2X1 U1130 ( .A(arr[548]), .B(n2766), .Y(n5074) );
  OAI21X1 U1131 ( .A(n4509), .B(n2767), .C(n5075), .Y(n7307) );
  NAND2X1 U1132 ( .A(arr[549]), .B(n2767), .Y(n5075) );
  OAI21X1 U1133 ( .A(n4511), .B(n2767), .C(n5076), .Y(n7308) );
  NAND2X1 U1134 ( .A(arr[550]), .B(n2768), .Y(n5076) );
  OAI21X1 U1135 ( .A(n4513), .B(n2766), .C(n5077), .Y(n7309) );
  NAND2X1 U1136 ( .A(arr[551]), .B(n2768), .Y(n5077) );
  OAI21X1 U1137 ( .A(n4515), .B(n2767), .C(n5078), .Y(n7310) );
  NAND2X1 U1138 ( .A(arr[552]), .B(n2768), .Y(n5078) );
  OAI21X1 U1139 ( .A(n4517), .B(n2766), .C(n5079), .Y(n7311) );
  NAND2X1 U1140 ( .A(arr[553]), .B(n2767), .Y(n5079) );
  OAI21X1 U1141 ( .A(n4519), .B(n2766), .C(n5080), .Y(n7312) );
  NAND2X1 U1142 ( .A(arr[554]), .B(n2766), .Y(n5080) );
  OAI21X1 U1143 ( .A(n4521), .B(n2766), .C(n5081), .Y(n7313) );
  NAND2X1 U1144 ( .A(arr[555]), .B(n2768), .Y(n5081) );
  OAI21X1 U1145 ( .A(n4523), .B(n2766), .C(n5082), .Y(n7314) );
  NAND2X1 U1146 ( .A(arr[556]), .B(n2767), .Y(n5082) );
  OAI21X1 U1147 ( .A(n4525), .B(n2766), .C(n5083), .Y(n7315) );
  NAND2X1 U1148 ( .A(arr[557]), .B(n2767), .Y(n5083) );
  OAI21X1 U1149 ( .A(n4527), .B(n2766), .C(n5084), .Y(n7316) );
  NAND2X1 U1150 ( .A(arr[558]), .B(n2766), .Y(n5084) );
  OAI21X1 U1151 ( .A(n4529), .B(n2766), .C(n5085), .Y(n7317) );
  NAND2X1 U1152 ( .A(arr[559]), .B(n2768), .Y(n5085) );
  OAI21X1 U1153 ( .A(n4531), .B(n2766), .C(n5086), .Y(n7318) );
  NAND2X1 U1154 ( .A(arr[560]), .B(n2766), .Y(n5086) );
  OAI21X1 U1156 ( .A(n4467), .B(n2765), .C(n5089), .Y(n7319) );
  NAND2X1 U1157 ( .A(arr[561]), .B(n2764), .Y(n5089) );
  OAI21X1 U1158 ( .A(n4469), .B(n2763), .C(n5090), .Y(n7320) );
  NAND2X1 U1159 ( .A(arr[562]), .B(n2764), .Y(n5090) );
  OAI21X1 U1160 ( .A(n4471), .B(n2763), .C(n5091), .Y(n7321) );
  NAND2X1 U1161 ( .A(arr[563]), .B(n2764), .Y(n5091) );
  OAI21X1 U1162 ( .A(n4473), .B(n2763), .C(n5092), .Y(n7322) );
  NAND2X1 U1163 ( .A(arr[564]), .B(n2764), .Y(n5092) );
  OAI21X1 U1164 ( .A(n4475), .B(n2763), .C(n5093), .Y(n7323) );
  NAND2X1 U1165 ( .A(arr[565]), .B(n2764), .Y(n5093) );
  OAI21X1 U1166 ( .A(n4477), .B(n2763), .C(n5094), .Y(n7324) );
  NAND2X1 U1167 ( .A(arr[566]), .B(n2765), .Y(n5094) );
  OAI21X1 U1168 ( .A(n4479), .B(n2763), .C(n5095), .Y(n7325) );
  NAND2X1 U1169 ( .A(arr[567]), .B(n2765), .Y(n5095) );
  OAI21X1 U1170 ( .A(n4481), .B(n2764), .C(n5096), .Y(n7326) );
  NAND2X1 U1171 ( .A(arr[568]), .B(n2764), .Y(n5096) );
  OAI21X1 U1172 ( .A(n4483), .B(n2763), .C(n5097), .Y(n7327) );
  NAND2X1 U1173 ( .A(arr[569]), .B(n2764), .Y(n5097) );
  OAI21X1 U1174 ( .A(n4485), .B(n2764), .C(n5098), .Y(n7328) );
  NAND2X1 U1175 ( .A(arr[570]), .B(n2765), .Y(n5098) );
  OAI21X1 U1176 ( .A(n4487), .B(n2764), .C(n5099), .Y(n7329) );
  NAND2X1 U1177 ( .A(arr[571]), .B(n2765), .Y(n5099) );
  OAI21X1 U1178 ( .A(n4489), .B(n2763), .C(n5100), .Y(n7330) );
  NAND2X1 U1179 ( .A(arr[572]), .B(n2765), .Y(n5100) );
  OAI21X1 U1180 ( .A(n4491), .B(n2764), .C(n5101), .Y(n7331) );
  NAND2X1 U1181 ( .A(arr[573]), .B(n2765), .Y(n5101) );
  OAI21X1 U1182 ( .A(n4493), .B(n2764), .C(n5102), .Y(n7332) );
  NAND2X1 U1183 ( .A(arr[574]), .B(n2765), .Y(n5102) );
  OAI21X1 U1184 ( .A(n4495), .B(n2763), .C(n5103), .Y(n7333) );
  NAND2X1 U1185 ( .A(arr[575]), .B(n2765), .Y(n5103) );
  OAI21X1 U1186 ( .A(n4497), .B(n2764), .C(n5104), .Y(n7334) );
  NAND2X1 U1187 ( .A(arr[576]), .B(n2765), .Y(n5104) );
  OAI21X1 U1188 ( .A(n4499), .B(n2764), .C(n5105), .Y(n7335) );
  NAND2X1 U1189 ( .A(arr[577]), .B(n2765), .Y(n5105) );
  OAI21X1 U1190 ( .A(n4501), .B(n2763), .C(n5106), .Y(n7336) );
  NAND2X1 U1191 ( .A(arr[578]), .B(n2765), .Y(n5106) );
  OAI21X1 U1192 ( .A(n4503), .B(n2763), .C(n5107), .Y(n7337) );
  NAND2X1 U1193 ( .A(arr[579]), .B(n2765), .Y(n5107) );
  OAI21X1 U1194 ( .A(n4505), .B(n2763), .C(n5108), .Y(n7338) );
  NAND2X1 U1195 ( .A(arr[580]), .B(n2765), .Y(n5108) );
  OAI21X1 U1196 ( .A(n4507), .B(n2763), .C(n5109), .Y(n7339) );
  NAND2X1 U1197 ( .A(arr[581]), .B(n2765), .Y(n5109) );
  OAI21X1 U1198 ( .A(n4509), .B(n2763), .C(n5110), .Y(n7340) );
  NAND2X1 U1199 ( .A(arr[582]), .B(n2765), .Y(n5110) );
  OAI21X1 U1200 ( .A(n4511), .B(n2763), .C(n5111), .Y(n7341) );
  NAND2X1 U1201 ( .A(arr[583]), .B(n2765), .Y(n5111) );
  OAI21X1 U1202 ( .A(n4513), .B(n2765), .C(n5112), .Y(n7342) );
  NAND2X1 U1203 ( .A(arr[584]), .B(n2765), .Y(n5112) );
  OAI21X1 U1204 ( .A(n4515), .B(n2763), .C(n5113), .Y(n7343) );
  NAND2X1 U1205 ( .A(arr[585]), .B(n2765), .Y(n5113) );
  OAI21X1 U1206 ( .A(n4517), .B(n2764), .C(n5114), .Y(n7344) );
  NAND2X1 U1207 ( .A(arr[586]), .B(n2765), .Y(n5114) );
  OAI21X1 U1208 ( .A(n4519), .B(n2763), .C(n5115), .Y(n7345) );
  NAND2X1 U1209 ( .A(arr[587]), .B(n2764), .Y(n5115) );
  OAI21X1 U1210 ( .A(n4521), .B(n2764), .C(n5116), .Y(n7346) );
  NAND2X1 U1211 ( .A(arr[588]), .B(n2765), .Y(n5116) );
  OAI21X1 U1212 ( .A(n4523), .B(n2763), .C(n5117), .Y(n7347) );
  NAND2X1 U1213 ( .A(arr[589]), .B(n2764), .Y(n5117) );
  OAI21X1 U1214 ( .A(n4525), .B(n2763), .C(n5118), .Y(n7348) );
  NAND2X1 U1215 ( .A(arr[590]), .B(n2765), .Y(n5118) );
  OAI21X1 U1216 ( .A(n4527), .B(n2763), .C(n5119), .Y(n7349) );
  NAND2X1 U1217 ( .A(arr[591]), .B(n2764), .Y(n5119) );
  OAI21X1 U1218 ( .A(n4529), .B(n2763), .C(n5120), .Y(n7350) );
  NAND2X1 U1219 ( .A(arr[592]), .B(n2764), .Y(n5120) );
  OAI21X1 U1220 ( .A(n4531), .B(n2763), .C(n5121), .Y(n7351) );
  NAND2X1 U1221 ( .A(arr[593]), .B(n2765), .Y(n5121) );
  OAI21X1 U1223 ( .A(n4467), .B(n2760), .C(n5123), .Y(n7352) );
  NAND2X1 U1224 ( .A(arr[594]), .B(n2762), .Y(n5123) );
  OAI21X1 U1225 ( .A(n4469), .B(n2760), .C(n5124), .Y(n7353) );
  NAND2X1 U1226 ( .A(arr[595]), .B(n2762), .Y(n5124) );
  OAI21X1 U1227 ( .A(n4471), .B(n2760), .C(n5125), .Y(n7354) );
  NAND2X1 U1228 ( .A(arr[596]), .B(n2762), .Y(n5125) );
  OAI21X1 U1229 ( .A(n4473), .B(n2760), .C(n5126), .Y(n7355) );
  NAND2X1 U1230 ( .A(arr[597]), .B(n2762), .Y(n5126) );
  OAI21X1 U1231 ( .A(n4475), .B(n2761), .C(n5127), .Y(n7356) );
  NAND2X1 U1232 ( .A(arr[598]), .B(n2762), .Y(n5127) );
  OAI21X1 U1233 ( .A(n4477), .B(n2761), .C(n5128), .Y(n7357) );
  NAND2X1 U1234 ( .A(arr[599]), .B(n2761), .Y(n5128) );
  OAI21X1 U1235 ( .A(n4479), .B(n2761), .C(n5129), .Y(n7358) );
  NAND2X1 U1236 ( .A(arr[600]), .B(n2762), .Y(n5129) );
  OAI21X1 U1237 ( .A(n4481), .B(n2762), .C(n5130), .Y(n7359) );
  NAND2X1 U1238 ( .A(arr[601]), .B(n2762), .Y(n5130) );
  OAI21X1 U1239 ( .A(n4483), .B(n2761), .C(n5131), .Y(n7360) );
  NAND2X1 U1240 ( .A(arr[602]), .B(n2762), .Y(n5131) );
  OAI21X1 U1241 ( .A(n4485), .B(n2762), .C(n5132), .Y(n7361) );
  NAND2X1 U1242 ( .A(arr[603]), .B(n2760), .Y(n5132) );
  OAI21X1 U1243 ( .A(n4487), .B(n2762), .C(n5133), .Y(n7362) );
  NAND2X1 U1244 ( .A(arr[604]), .B(n2762), .Y(n5133) );
  OAI21X1 U1245 ( .A(n4489), .B(n2761), .C(n5134), .Y(n7363) );
  NAND2X1 U1246 ( .A(arr[605]), .B(n2760), .Y(n5134) );
  OAI21X1 U1247 ( .A(n4491), .B(n2762), .C(n5135), .Y(n7364) );
  NAND2X1 U1248 ( .A(arr[606]), .B(n2761), .Y(n5135) );
  OAI21X1 U1249 ( .A(n4493), .B(n2762), .C(n5136), .Y(n7365) );
  NAND2X1 U1250 ( .A(arr[607]), .B(n2761), .Y(n5136) );
  OAI21X1 U1251 ( .A(n4495), .B(n2761), .C(n5137), .Y(n7366) );
  NAND2X1 U1252 ( .A(arr[608]), .B(n2762), .Y(n5137) );
  OAI21X1 U1253 ( .A(n4497), .B(n2762), .C(n5138), .Y(n7367) );
  NAND2X1 U1254 ( .A(arr[609]), .B(n2760), .Y(n5138) );
  OAI21X1 U1255 ( .A(n4499), .B(n2762), .C(n5139), .Y(n7368) );
  NAND2X1 U1256 ( .A(arr[610]), .B(n2762), .Y(n5139) );
  OAI21X1 U1257 ( .A(n4501), .B(n2761), .C(n5140), .Y(n7369) );
  NAND2X1 U1258 ( .A(arr[611]), .B(n2760), .Y(n5140) );
  OAI21X1 U1259 ( .A(n4503), .B(n2761), .C(n5141), .Y(n7370) );
  NAND2X1 U1260 ( .A(arr[612]), .B(n2761), .Y(n5141) );
  OAI21X1 U1261 ( .A(n4505), .B(n2761), .C(n5142), .Y(n7371) );
  NAND2X1 U1262 ( .A(arr[613]), .B(n2762), .Y(n5142) );
  OAI21X1 U1263 ( .A(n4507), .B(n2761), .C(n5143), .Y(n7372) );
  NAND2X1 U1264 ( .A(arr[614]), .B(n2760), .Y(n5143) );
  OAI21X1 U1265 ( .A(n4509), .B(n2761), .C(n5144), .Y(n7373) );
  NAND2X1 U1266 ( .A(arr[615]), .B(n2761), .Y(n5144) );
  OAI21X1 U1267 ( .A(n4511), .B(n2761), .C(n5145), .Y(n7374) );
  NAND2X1 U1268 ( .A(arr[616]), .B(n2762), .Y(n5145) );
  OAI21X1 U1269 ( .A(n4513), .B(n2760), .C(n5146), .Y(n7375) );
  NAND2X1 U1270 ( .A(arr[617]), .B(n2762), .Y(n5146) );
  OAI21X1 U1271 ( .A(n4515), .B(n2761), .C(n5147), .Y(n7376) );
  NAND2X1 U1272 ( .A(arr[618]), .B(n2762), .Y(n5147) );
  OAI21X1 U1273 ( .A(n4517), .B(n2760), .C(n5148), .Y(n7377) );
  NAND2X1 U1274 ( .A(arr[619]), .B(n2761), .Y(n5148) );
  OAI21X1 U1275 ( .A(n4519), .B(n2760), .C(n5149), .Y(n7378) );
  NAND2X1 U1276 ( .A(arr[620]), .B(n2760), .Y(n5149) );
  OAI21X1 U1277 ( .A(n4521), .B(n2760), .C(n5150), .Y(n7379) );
  NAND2X1 U1278 ( .A(arr[621]), .B(n2762), .Y(n5150) );
  OAI21X1 U1279 ( .A(n4523), .B(n2760), .C(n5151), .Y(n7380) );
  NAND2X1 U1280 ( .A(arr[622]), .B(n2761), .Y(n5151) );
  OAI21X1 U1281 ( .A(n4525), .B(n2760), .C(n5152), .Y(n7381) );
  NAND2X1 U1282 ( .A(arr[623]), .B(n2761), .Y(n5152) );
  OAI21X1 U1283 ( .A(n4527), .B(n2760), .C(n5153), .Y(n7382) );
  NAND2X1 U1284 ( .A(arr[624]), .B(n2760), .Y(n5153) );
  OAI21X1 U1285 ( .A(n4529), .B(n2760), .C(n5154), .Y(n7383) );
  NAND2X1 U1286 ( .A(arr[625]), .B(n2762), .Y(n5154) );
  OAI21X1 U1287 ( .A(n4531), .B(n2760), .C(n5155), .Y(n7384) );
  NAND2X1 U1288 ( .A(arr[626]), .B(n2760), .Y(n5155) );
  OAI21X1 U1290 ( .A(n4467), .B(n2759), .C(n5158), .Y(n7385) );
  NAND2X1 U1291 ( .A(arr[627]), .B(n2758), .Y(n5158) );
  OAI21X1 U1292 ( .A(n4469), .B(n2757), .C(n5159), .Y(n7386) );
  NAND2X1 U1293 ( .A(arr[628]), .B(n2758), .Y(n5159) );
  OAI21X1 U1294 ( .A(n4471), .B(n2757), .C(n5160), .Y(n7387) );
  NAND2X1 U1295 ( .A(arr[629]), .B(n2758), .Y(n5160) );
  OAI21X1 U1296 ( .A(n4473), .B(n2757), .C(n5161), .Y(n7388) );
  NAND2X1 U1297 ( .A(arr[630]), .B(n2758), .Y(n5161) );
  OAI21X1 U1298 ( .A(n4475), .B(n2757), .C(n5162), .Y(n7389) );
  NAND2X1 U1299 ( .A(arr[631]), .B(n2758), .Y(n5162) );
  OAI21X1 U1300 ( .A(n4477), .B(n2757), .C(n5163), .Y(n7390) );
  NAND2X1 U1301 ( .A(arr[632]), .B(n2759), .Y(n5163) );
  OAI21X1 U1302 ( .A(n4479), .B(n2757), .C(n5164), .Y(n7391) );
  NAND2X1 U1303 ( .A(arr[633]), .B(n2759), .Y(n5164) );
  OAI21X1 U1304 ( .A(n4481), .B(n2758), .C(n5165), .Y(n7392) );
  NAND2X1 U1305 ( .A(arr[634]), .B(n2758), .Y(n5165) );
  OAI21X1 U1306 ( .A(n4483), .B(n2757), .C(n5166), .Y(n7393) );
  NAND2X1 U1307 ( .A(arr[635]), .B(n2758), .Y(n5166) );
  OAI21X1 U1308 ( .A(n4485), .B(n2758), .C(n5167), .Y(n7394) );
  NAND2X1 U1309 ( .A(arr[636]), .B(n2759), .Y(n5167) );
  OAI21X1 U1310 ( .A(n4487), .B(n2758), .C(n5168), .Y(n7395) );
  NAND2X1 U1311 ( .A(arr[637]), .B(n2759), .Y(n5168) );
  OAI21X1 U1312 ( .A(n4489), .B(n2757), .C(n5169), .Y(n7396) );
  NAND2X1 U1313 ( .A(arr[638]), .B(n2759), .Y(n5169) );
  OAI21X1 U1314 ( .A(n4491), .B(n2758), .C(n5170), .Y(n7397) );
  NAND2X1 U1315 ( .A(arr[639]), .B(n2759), .Y(n5170) );
  OAI21X1 U1316 ( .A(n4493), .B(n2758), .C(n5171), .Y(n7398) );
  NAND2X1 U1317 ( .A(arr[640]), .B(n2759), .Y(n5171) );
  OAI21X1 U1318 ( .A(n4495), .B(n2757), .C(n5172), .Y(n7399) );
  NAND2X1 U1319 ( .A(arr[641]), .B(n2759), .Y(n5172) );
  OAI21X1 U1320 ( .A(n4497), .B(n2758), .C(n5173), .Y(n7400) );
  NAND2X1 U1321 ( .A(arr[642]), .B(n2759), .Y(n5173) );
  OAI21X1 U1322 ( .A(n4499), .B(n2758), .C(n5174), .Y(n7401) );
  NAND2X1 U1323 ( .A(arr[643]), .B(n2759), .Y(n5174) );
  OAI21X1 U1324 ( .A(n4501), .B(n2757), .C(n5175), .Y(n7402) );
  NAND2X1 U1325 ( .A(arr[644]), .B(n2759), .Y(n5175) );
  OAI21X1 U1326 ( .A(n4503), .B(n2757), .C(n5176), .Y(n7403) );
  NAND2X1 U1327 ( .A(arr[645]), .B(n2759), .Y(n5176) );
  OAI21X1 U1328 ( .A(n4505), .B(n2757), .C(n5177), .Y(n7404) );
  NAND2X1 U1329 ( .A(arr[646]), .B(n2759), .Y(n5177) );
  OAI21X1 U1330 ( .A(n4507), .B(n2757), .C(n5178), .Y(n7405) );
  NAND2X1 U1331 ( .A(arr[647]), .B(n2759), .Y(n5178) );
  OAI21X1 U1332 ( .A(n4509), .B(n2757), .C(n5179), .Y(n7406) );
  NAND2X1 U1333 ( .A(arr[648]), .B(n2759), .Y(n5179) );
  OAI21X1 U1334 ( .A(n4511), .B(n2757), .C(n5180), .Y(n7407) );
  NAND2X1 U1335 ( .A(arr[649]), .B(n2759), .Y(n5180) );
  OAI21X1 U1336 ( .A(n4513), .B(n2759), .C(n5181), .Y(n7408) );
  NAND2X1 U1337 ( .A(arr[650]), .B(n2759), .Y(n5181) );
  OAI21X1 U1338 ( .A(n4515), .B(n2757), .C(n5182), .Y(n7409) );
  NAND2X1 U1339 ( .A(arr[651]), .B(n2759), .Y(n5182) );
  OAI21X1 U1340 ( .A(n4517), .B(n2758), .C(n5183), .Y(n7410) );
  NAND2X1 U1341 ( .A(arr[652]), .B(n2759), .Y(n5183) );
  OAI21X1 U1342 ( .A(n4519), .B(n2757), .C(n5184), .Y(n7411) );
  NAND2X1 U1343 ( .A(arr[653]), .B(n2758), .Y(n5184) );
  OAI21X1 U1344 ( .A(n4521), .B(n2758), .C(n5185), .Y(n7412) );
  NAND2X1 U1345 ( .A(arr[654]), .B(n2759), .Y(n5185) );
  OAI21X1 U1346 ( .A(n4523), .B(n2757), .C(n5186), .Y(n7413) );
  NAND2X1 U1347 ( .A(arr[655]), .B(n2758), .Y(n5186) );
  OAI21X1 U1348 ( .A(n4525), .B(n2757), .C(n5187), .Y(n7414) );
  NAND2X1 U1349 ( .A(arr[656]), .B(n2759), .Y(n5187) );
  OAI21X1 U1350 ( .A(n4527), .B(n2757), .C(n5188), .Y(n7415) );
  NAND2X1 U1351 ( .A(arr[657]), .B(n2758), .Y(n5188) );
  OAI21X1 U1352 ( .A(n4529), .B(n2757), .C(n5189), .Y(n7416) );
  NAND2X1 U1353 ( .A(arr[658]), .B(n2758), .Y(n5189) );
  OAI21X1 U1354 ( .A(n4531), .B(n2757), .C(n5190), .Y(n7417) );
  NAND2X1 U1355 ( .A(arr[659]), .B(n2759), .Y(n5190) );
  OAI21X1 U1357 ( .A(n4467), .B(n2754), .C(n5192), .Y(n7418) );
  NAND2X1 U1358 ( .A(arr[660]), .B(n2756), .Y(n5192) );
  OAI21X1 U1359 ( .A(n4469), .B(n2754), .C(n5193), .Y(n7419) );
  NAND2X1 U1360 ( .A(arr[661]), .B(n2756), .Y(n5193) );
  OAI21X1 U1361 ( .A(n4471), .B(n2754), .C(n5194), .Y(n7420) );
  NAND2X1 U1362 ( .A(arr[662]), .B(n2756), .Y(n5194) );
  OAI21X1 U1363 ( .A(n4473), .B(n2754), .C(n5195), .Y(n7421) );
  NAND2X1 U1364 ( .A(arr[663]), .B(n2756), .Y(n5195) );
  OAI21X1 U1365 ( .A(n4475), .B(n2755), .C(n5196), .Y(n7422) );
  NAND2X1 U1366 ( .A(arr[664]), .B(n2756), .Y(n5196) );
  OAI21X1 U1367 ( .A(n4477), .B(n2755), .C(n5197), .Y(n7423) );
  NAND2X1 U1368 ( .A(arr[665]), .B(n2755), .Y(n5197) );
  OAI21X1 U1369 ( .A(n4479), .B(n2755), .C(n5198), .Y(n7424) );
  NAND2X1 U1370 ( .A(arr[666]), .B(n2756), .Y(n5198) );
  OAI21X1 U1371 ( .A(n4481), .B(n2756), .C(n5199), .Y(n7425) );
  NAND2X1 U1372 ( .A(arr[667]), .B(n2756), .Y(n5199) );
  OAI21X1 U1373 ( .A(n4483), .B(n2755), .C(n5200), .Y(n7426) );
  NAND2X1 U1374 ( .A(arr[668]), .B(n2756), .Y(n5200) );
  OAI21X1 U1375 ( .A(n4485), .B(n2756), .C(n5201), .Y(n7427) );
  NAND2X1 U1376 ( .A(arr[669]), .B(n2754), .Y(n5201) );
  OAI21X1 U1377 ( .A(n4487), .B(n2756), .C(n5202), .Y(n7428) );
  NAND2X1 U1378 ( .A(arr[670]), .B(n2756), .Y(n5202) );
  OAI21X1 U1379 ( .A(n4489), .B(n2755), .C(n5203), .Y(n7429) );
  NAND2X1 U1380 ( .A(arr[671]), .B(n2754), .Y(n5203) );
  OAI21X1 U1381 ( .A(n4491), .B(n2756), .C(n5204), .Y(n7430) );
  NAND2X1 U1382 ( .A(arr[672]), .B(n2755), .Y(n5204) );
  OAI21X1 U1383 ( .A(n4493), .B(n2756), .C(n5205), .Y(n7431) );
  NAND2X1 U1384 ( .A(arr[673]), .B(n2755), .Y(n5205) );
  OAI21X1 U1385 ( .A(n4495), .B(n2755), .C(n5206), .Y(n7432) );
  NAND2X1 U1386 ( .A(arr[674]), .B(n2756), .Y(n5206) );
  OAI21X1 U1387 ( .A(n4497), .B(n2756), .C(n5207), .Y(n7433) );
  NAND2X1 U1388 ( .A(arr[675]), .B(n2754), .Y(n5207) );
  OAI21X1 U1389 ( .A(n4499), .B(n2756), .C(n5208), .Y(n7434) );
  NAND2X1 U1390 ( .A(arr[676]), .B(n2756), .Y(n5208) );
  OAI21X1 U1391 ( .A(n4501), .B(n2755), .C(n5209), .Y(n7435) );
  NAND2X1 U1392 ( .A(arr[677]), .B(n2754), .Y(n5209) );
  OAI21X1 U1393 ( .A(n4503), .B(n2755), .C(n5210), .Y(n7436) );
  NAND2X1 U1394 ( .A(arr[678]), .B(n2755), .Y(n5210) );
  OAI21X1 U1395 ( .A(n4505), .B(n2755), .C(n5211), .Y(n7437) );
  NAND2X1 U1396 ( .A(arr[679]), .B(n2756), .Y(n5211) );
  OAI21X1 U1397 ( .A(n4507), .B(n2755), .C(n5212), .Y(n7438) );
  NAND2X1 U1398 ( .A(arr[680]), .B(n2754), .Y(n5212) );
  OAI21X1 U1399 ( .A(n4509), .B(n2755), .C(n5213), .Y(n7439) );
  NAND2X1 U1400 ( .A(arr[681]), .B(n2755), .Y(n5213) );
  OAI21X1 U1401 ( .A(n4511), .B(n2755), .C(n5214), .Y(n7440) );
  NAND2X1 U1402 ( .A(arr[682]), .B(n2756), .Y(n5214) );
  OAI21X1 U1403 ( .A(n4513), .B(n2754), .C(n5215), .Y(n7441) );
  NAND2X1 U1404 ( .A(arr[683]), .B(n2756), .Y(n5215) );
  OAI21X1 U1405 ( .A(n4515), .B(n2755), .C(n5216), .Y(n7442) );
  NAND2X1 U1406 ( .A(arr[684]), .B(n2756), .Y(n5216) );
  OAI21X1 U1407 ( .A(n4517), .B(n2754), .C(n5217), .Y(n7443) );
  NAND2X1 U1408 ( .A(arr[685]), .B(n2755), .Y(n5217) );
  OAI21X1 U1409 ( .A(n4519), .B(n2754), .C(n5218), .Y(n7444) );
  NAND2X1 U1410 ( .A(arr[686]), .B(n2754), .Y(n5218) );
  OAI21X1 U1411 ( .A(n4521), .B(n2754), .C(n5219), .Y(n7445) );
  NAND2X1 U1412 ( .A(arr[687]), .B(n2756), .Y(n5219) );
  OAI21X1 U1413 ( .A(n4523), .B(n2754), .C(n5220), .Y(n7446) );
  NAND2X1 U1414 ( .A(arr[688]), .B(n2755), .Y(n5220) );
  OAI21X1 U1415 ( .A(n4525), .B(n2754), .C(n5221), .Y(n7447) );
  NAND2X1 U1416 ( .A(arr[689]), .B(n2755), .Y(n5221) );
  OAI21X1 U1417 ( .A(n4527), .B(n2754), .C(n5222), .Y(n7448) );
  NAND2X1 U1418 ( .A(arr[690]), .B(n2754), .Y(n5222) );
  OAI21X1 U1419 ( .A(n4529), .B(n2754), .C(n5223), .Y(n7449) );
  NAND2X1 U1420 ( .A(arr[691]), .B(n2756), .Y(n5223) );
  OAI21X1 U1421 ( .A(n4531), .B(n2754), .C(n5224), .Y(n7450) );
  NAND2X1 U1422 ( .A(arr[692]), .B(n2754), .Y(n5224) );
  OAI21X1 U1424 ( .A(n4467), .B(n2753), .C(n5227), .Y(n7451) );
  NAND2X1 U1425 ( .A(arr[693]), .B(n2752), .Y(n5227) );
  OAI21X1 U1426 ( .A(n4469), .B(n2751), .C(n5228), .Y(n7452) );
  NAND2X1 U1427 ( .A(arr[694]), .B(n2752), .Y(n5228) );
  OAI21X1 U1428 ( .A(n4471), .B(n2751), .C(n5229), .Y(n7453) );
  NAND2X1 U1429 ( .A(arr[695]), .B(n2752), .Y(n5229) );
  OAI21X1 U1430 ( .A(n4473), .B(n2751), .C(n5230), .Y(n7454) );
  NAND2X1 U1431 ( .A(arr[696]), .B(n2752), .Y(n5230) );
  OAI21X1 U1432 ( .A(n4475), .B(n2751), .C(n5231), .Y(n7455) );
  NAND2X1 U1433 ( .A(arr[697]), .B(n2752), .Y(n5231) );
  OAI21X1 U1434 ( .A(n4477), .B(n2751), .C(n5232), .Y(n7456) );
  NAND2X1 U1435 ( .A(arr[698]), .B(n2753), .Y(n5232) );
  OAI21X1 U1436 ( .A(n4479), .B(n2751), .C(n5233), .Y(n7457) );
  NAND2X1 U1437 ( .A(arr[699]), .B(n2753), .Y(n5233) );
  OAI21X1 U1438 ( .A(n4481), .B(n2752), .C(n5234), .Y(n7458) );
  NAND2X1 U1439 ( .A(arr[700]), .B(n2752), .Y(n5234) );
  OAI21X1 U1440 ( .A(n4483), .B(n2751), .C(n5235), .Y(n7459) );
  NAND2X1 U1441 ( .A(arr[701]), .B(n2752), .Y(n5235) );
  OAI21X1 U1442 ( .A(n4485), .B(n2752), .C(n5236), .Y(n7460) );
  NAND2X1 U1443 ( .A(arr[702]), .B(n2753), .Y(n5236) );
  OAI21X1 U1444 ( .A(n4487), .B(n2752), .C(n5237), .Y(n7461) );
  NAND2X1 U1445 ( .A(arr[703]), .B(n2753), .Y(n5237) );
  OAI21X1 U1446 ( .A(n4489), .B(n2751), .C(n5238), .Y(n7462) );
  NAND2X1 U1447 ( .A(arr[704]), .B(n2753), .Y(n5238) );
  OAI21X1 U1448 ( .A(n4491), .B(n2752), .C(n5239), .Y(n7463) );
  NAND2X1 U1449 ( .A(arr[705]), .B(n2753), .Y(n5239) );
  OAI21X1 U1450 ( .A(n4493), .B(n2752), .C(n5240), .Y(n7464) );
  NAND2X1 U1451 ( .A(arr[706]), .B(n2753), .Y(n5240) );
  OAI21X1 U1452 ( .A(n4495), .B(n2751), .C(n5241), .Y(n7465) );
  NAND2X1 U1453 ( .A(arr[707]), .B(n2753), .Y(n5241) );
  OAI21X1 U1454 ( .A(n4497), .B(n2752), .C(n5242), .Y(n7466) );
  NAND2X1 U1455 ( .A(arr[708]), .B(n2753), .Y(n5242) );
  OAI21X1 U1456 ( .A(n4499), .B(n2752), .C(n5243), .Y(n7467) );
  NAND2X1 U1457 ( .A(arr[709]), .B(n2753), .Y(n5243) );
  OAI21X1 U1458 ( .A(n4501), .B(n2751), .C(n5244), .Y(n7468) );
  NAND2X1 U1459 ( .A(arr[710]), .B(n2753), .Y(n5244) );
  OAI21X1 U1460 ( .A(n4503), .B(n2751), .C(n5245), .Y(n7469) );
  NAND2X1 U1461 ( .A(arr[711]), .B(n2753), .Y(n5245) );
  OAI21X1 U1462 ( .A(n4505), .B(n2751), .C(n5246), .Y(n7470) );
  NAND2X1 U1463 ( .A(arr[712]), .B(n2753), .Y(n5246) );
  OAI21X1 U1464 ( .A(n4507), .B(n2751), .C(n5247), .Y(n7471) );
  NAND2X1 U1465 ( .A(arr[713]), .B(n2753), .Y(n5247) );
  OAI21X1 U1466 ( .A(n4509), .B(n2751), .C(n5248), .Y(n7472) );
  NAND2X1 U1467 ( .A(arr[714]), .B(n2753), .Y(n5248) );
  OAI21X1 U1468 ( .A(n4511), .B(n2751), .C(n5249), .Y(n7473) );
  NAND2X1 U1469 ( .A(arr[715]), .B(n2753), .Y(n5249) );
  OAI21X1 U1470 ( .A(n4513), .B(n2753), .C(n5250), .Y(n7474) );
  NAND2X1 U1471 ( .A(arr[716]), .B(n2753), .Y(n5250) );
  OAI21X1 U1472 ( .A(n4515), .B(n2751), .C(n5251), .Y(n7475) );
  NAND2X1 U1473 ( .A(arr[717]), .B(n2753), .Y(n5251) );
  OAI21X1 U1474 ( .A(n4517), .B(n2752), .C(n5252), .Y(n7476) );
  NAND2X1 U1475 ( .A(arr[718]), .B(n2753), .Y(n5252) );
  OAI21X1 U1476 ( .A(n4519), .B(n2751), .C(n5253), .Y(n7477) );
  NAND2X1 U1477 ( .A(arr[719]), .B(n2752), .Y(n5253) );
  OAI21X1 U1478 ( .A(n4521), .B(n2752), .C(n5254), .Y(n7478) );
  NAND2X1 U1479 ( .A(arr[720]), .B(n2753), .Y(n5254) );
  OAI21X1 U1480 ( .A(n4523), .B(n2751), .C(n5255), .Y(n7479) );
  NAND2X1 U1481 ( .A(arr[721]), .B(n2752), .Y(n5255) );
  OAI21X1 U1482 ( .A(n4525), .B(n2751), .C(n5256), .Y(n7480) );
  NAND2X1 U1483 ( .A(arr[722]), .B(n2753), .Y(n5256) );
  OAI21X1 U1484 ( .A(n4527), .B(n2751), .C(n5257), .Y(n7481) );
  NAND2X1 U1485 ( .A(arr[723]), .B(n2752), .Y(n5257) );
  OAI21X1 U1486 ( .A(n4529), .B(n2751), .C(n5258), .Y(n7482) );
  NAND2X1 U1487 ( .A(arr[724]), .B(n2752), .Y(n5258) );
  OAI21X1 U1488 ( .A(n4531), .B(n2751), .C(n5259), .Y(n7483) );
  NAND2X1 U1489 ( .A(arr[725]), .B(n2753), .Y(n5259) );
  OAI21X1 U1491 ( .A(n4467), .B(n2748), .C(n5261), .Y(n7484) );
  NAND2X1 U1492 ( .A(arr[726]), .B(n2750), .Y(n5261) );
  OAI21X1 U1493 ( .A(n4469), .B(n2748), .C(n5262), .Y(n7485) );
  NAND2X1 U1494 ( .A(arr[727]), .B(n2750), .Y(n5262) );
  OAI21X1 U1495 ( .A(n4471), .B(n2748), .C(n5263), .Y(n7486) );
  NAND2X1 U1496 ( .A(arr[728]), .B(n2750), .Y(n5263) );
  OAI21X1 U1497 ( .A(n4473), .B(n2748), .C(n5264), .Y(n7487) );
  NAND2X1 U1498 ( .A(arr[729]), .B(n2750), .Y(n5264) );
  OAI21X1 U1499 ( .A(n4475), .B(n2749), .C(n5265), .Y(n7488) );
  NAND2X1 U1500 ( .A(arr[730]), .B(n2750), .Y(n5265) );
  OAI21X1 U1501 ( .A(n4477), .B(n2749), .C(n5266), .Y(n7489) );
  NAND2X1 U1502 ( .A(arr[731]), .B(n2749), .Y(n5266) );
  OAI21X1 U1503 ( .A(n4479), .B(n2749), .C(n5267), .Y(n7490) );
  NAND2X1 U1504 ( .A(arr[732]), .B(n2750), .Y(n5267) );
  OAI21X1 U1505 ( .A(n4481), .B(n2750), .C(n5268), .Y(n7491) );
  NAND2X1 U1506 ( .A(arr[733]), .B(n2750), .Y(n5268) );
  OAI21X1 U1507 ( .A(n4483), .B(n2749), .C(n5269), .Y(n7492) );
  NAND2X1 U1508 ( .A(arr[734]), .B(n2750), .Y(n5269) );
  OAI21X1 U1509 ( .A(n4485), .B(n2750), .C(n5270), .Y(n7493) );
  NAND2X1 U1510 ( .A(arr[735]), .B(n2748), .Y(n5270) );
  OAI21X1 U1511 ( .A(n4487), .B(n2750), .C(n5271), .Y(n7494) );
  NAND2X1 U1512 ( .A(arr[736]), .B(n2750), .Y(n5271) );
  OAI21X1 U1513 ( .A(n4489), .B(n2749), .C(n5272), .Y(n7495) );
  NAND2X1 U1514 ( .A(arr[737]), .B(n2748), .Y(n5272) );
  OAI21X1 U1515 ( .A(n4491), .B(n2750), .C(n5273), .Y(n7496) );
  NAND2X1 U1516 ( .A(arr[738]), .B(n2749), .Y(n5273) );
  OAI21X1 U1517 ( .A(n4493), .B(n2750), .C(n5274), .Y(n7497) );
  NAND2X1 U1518 ( .A(arr[739]), .B(n2749), .Y(n5274) );
  OAI21X1 U1519 ( .A(n4495), .B(n2749), .C(n5275), .Y(n7498) );
  NAND2X1 U1520 ( .A(arr[740]), .B(n2750), .Y(n5275) );
  OAI21X1 U1521 ( .A(n4497), .B(n2750), .C(n5276), .Y(n7499) );
  NAND2X1 U1522 ( .A(arr[741]), .B(n2748), .Y(n5276) );
  OAI21X1 U1523 ( .A(n4499), .B(n2750), .C(n5277), .Y(n7500) );
  NAND2X1 U1524 ( .A(arr[742]), .B(n2750), .Y(n5277) );
  OAI21X1 U1525 ( .A(n4501), .B(n2749), .C(n5278), .Y(n7501) );
  NAND2X1 U1526 ( .A(arr[743]), .B(n2748), .Y(n5278) );
  OAI21X1 U1527 ( .A(n4503), .B(n2749), .C(n5279), .Y(n7502) );
  NAND2X1 U1528 ( .A(arr[744]), .B(n2749), .Y(n5279) );
  OAI21X1 U1529 ( .A(n4505), .B(n2749), .C(n5280), .Y(n7503) );
  NAND2X1 U1530 ( .A(arr[745]), .B(n2750), .Y(n5280) );
  OAI21X1 U1531 ( .A(n4507), .B(n2749), .C(n5281), .Y(n7504) );
  NAND2X1 U1532 ( .A(arr[746]), .B(n2748), .Y(n5281) );
  OAI21X1 U1533 ( .A(n4509), .B(n2749), .C(n5282), .Y(n7505) );
  NAND2X1 U1534 ( .A(arr[747]), .B(n2749), .Y(n5282) );
  OAI21X1 U1535 ( .A(n4511), .B(n2749), .C(n5283), .Y(n7506) );
  NAND2X1 U1536 ( .A(arr[748]), .B(n2750), .Y(n5283) );
  OAI21X1 U1537 ( .A(n4513), .B(n2748), .C(n5284), .Y(n7507) );
  NAND2X1 U1538 ( .A(arr[749]), .B(n2750), .Y(n5284) );
  OAI21X1 U1539 ( .A(n4515), .B(n2749), .C(n5285), .Y(n7508) );
  NAND2X1 U1540 ( .A(arr[750]), .B(n2750), .Y(n5285) );
  OAI21X1 U1541 ( .A(n4517), .B(n2748), .C(n5286), .Y(n7509) );
  NAND2X1 U1542 ( .A(arr[751]), .B(n2749), .Y(n5286) );
  OAI21X1 U1543 ( .A(n4519), .B(n2748), .C(n5287), .Y(n7510) );
  NAND2X1 U1544 ( .A(arr[752]), .B(n2748), .Y(n5287) );
  OAI21X1 U1545 ( .A(n4521), .B(n2748), .C(n5288), .Y(n7511) );
  NAND2X1 U1546 ( .A(arr[753]), .B(n2750), .Y(n5288) );
  OAI21X1 U1547 ( .A(n4523), .B(n2748), .C(n5289), .Y(n7512) );
  NAND2X1 U1548 ( .A(arr[754]), .B(n2749), .Y(n5289) );
  OAI21X1 U1549 ( .A(n4525), .B(n2748), .C(n5290), .Y(n7513) );
  NAND2X1 U1550 ( .A(arr[755]), .B(n2749), .Y(n5290) );
  OAI21X1 U1551 ( .A(n4527), .B(n2748), .C(n5291), .Y(n7514) );
  NAND2X1 U1552 ( .A(arr[756]), .B(n2748), .Y(n5291) );
  OAI21X1 U1553 ( .A(n4529), .B(n2748), .C(n5292), .Y(n7515) );
  NAND2X1 U1554 ( .A(arr[757]), .B(n2750), .Y(n5292) );
  OAI21X1 U1555 ( .A(n4531), .B(n2748), .C(n5293), .Y(n7516) );
  NAND2X1 U1556 ( .A(arr[758]), .B(n2748), .Y(n5293) );
  OAI21X1 U1558 ( .A(n4467), .B(n2747), .C(n5296), .Y(n7517) );
  NAND2X1 U1559 ( .A(arr[759]), .B(n2746), .Y(n5296) );
  OAI21X1 U1560 ( .A(n4469), .B(n2745), .C(n5297), .Y(n7518) );
  NAND2X1 U1561 ( .A(arr[760]), .B(n2746), .Y(n5297) );
  OAI21X1 U1562 ( .A(n4471), .B(n2745), .C(n5298), .Y(n7519) );
  NAND2X1 U1563 ( .A(arr[761]), .B(n2746), .Y(n5298) );
  OAI21X1 U1564 ( .A(n4473), .B(n2745), .C(n5299), .Y(n7520) );
  NAND2X1 U1565 ( .A(arr[762]), .B(n2746), .Y(n5299) );
  OAI21X1 U1566 ( .A(n4475), .B(n2745), .C(n5300), .Y(n7521) );
  NAND2X1 U1567 ( .A(arr[763]), .B(n2746), .Y(n5300) );
  OAI21X1 U1568 ( .A(n4477), .B(n2745), .C(n5301), .Y(n7522) );
  NAND2X1 U1569 ( .A(arr[764]), .B(n2747), .Y(n5301) );
  OAI21X1 U1570 ( .A(n4479), .B(n2745), .C(n5302), .Y(n7523) );
  NAND2X1 U1571 ( .A(arr[765]), .B(n2747), .Y(n5302) );
  OAI21X1 U1572 ( .A(n4481), .B(n2746), .C(n5303), .Y(n7524) );
  NAND2X1 U1573 ( .A(arr[766]), .B(n2746), .Y(n5303) );
  OAI21X1 U1574 ( .A(n4483), .B(n2745), .C(n5304), .Y(n7525) );
  NAND2X1 U1575 ( .A(arr[767]), .B(n2746), .Y(n5304) );
  OAI21X1 U1576 ( .A(n4485), .B(n2746), .C(n5305), .Y(n7526) );
  NAND2X1 U1577 ( .A(arr[768]), .B(n2747), .Y(n5305) );
  OAI21X1 U1578 ( .A(n4487), .B(n2746), .C(n5306), .Y(n7527) );
  NAND2X1 U1579 ( .A(arr[769]), .B(n2747), .Y(n5306) );
  OAI21X1 U1580 ( .A(n4489), .B(n2745), .C(n5307), .Y(n7528) );
  NAND2X1 U1581 ( .A(arr[770]), .B(n2747), .Y(n5307) );
  OAI21X1 U1582 ( .A(n4491), .B(n2746), .C(n5308), .Y(n7529) );
  NAND2X1 U1583 ( .A(arr[771]), .B(n2747), .Y(n5308) );
  OAI21X1 U1584 ( .A(n4493), .B(n2746), .C(n5309), .Y(n7530) );
  NAND2X1 U1585 ( .A(arr[772]), .B(n2747), .Y(n5309) );
  OAI21X1 U1586 ( .A(n4495), .B(n2745), .C(n5310), .Y(n7531) );
  NAND2X1 U1587 ( .A(arr[773]), .B(n2747), .Y(n5310) );
  OAI21X1 U1588 ( .A(n4497), .B(n2746), .C(n5311), .Y(n7532) );
  NAND2X1 U1589 ( .A(arr[774]), .B(n2747), .Y(n5311) );
  OAI21X1 U1590 ( .A(n4499), .B(n2746), .C(n5312), .Y(n7533) );
  NAND2X1 U1591 ( .A(arr[775]), .B(n2747), .Y(n5312) );
  OAI21X1 U1592 ( .A(n4501), .B(n2745), .C(n5313), .Y(n7534) );
  NAND2X1 U1593 ( .A(arr[776]), .B(n2747), .Y(n5313) );
  OAI21X1 U1594 ( .A(n4503), .B(n2745), .C(n5314), .Y(n7535) );
  NAND2X1 U1595 ( .A(arr[777]), .B(n2747), .Y(n5314) );
  OAI21X1 U1596 ( .A(n4505), .B(n2745), .C(n5315), .Y(n7536) );
  NAND2X1 U1597 ( .A(arr[778]), .B(n2747), .Y(n5315) );
  OAI21X1 U1598 ( .A(n4507), .B(n2745), .C(n5316), .Y(n7537) );
  NAND2X1 U1599 ( .A(arr[779]), .B(n2747), .Y(n5316) );
  OAI21X1 U1600 ( .A(n4509), .B(n2745), .C(n5317), .Y(n7538) );
  NAND2X1 U1601 ( .A(arr[780]), .B(n2747), .Y(n5317) );
  OAI21X1 U1602 ( .A(n4511), .B(n2745), .C(n5318), .Y(n7539) );
  NAND2X1 U1603 ( .A(arr[781]), .B(n2747), .Y(n5318) );
  OAI21X1 U1604 ( .A(n4513), .B(n2747), .C(n5319), .Y(n7540) );
  NAND2X1 U1605 ( .A(arr[782]), .B(n2747), .Y(n5319) );
  OAI21X1 U1606 ( .A(n4515), .B(n2745), .C(n5320), .Y(n7541) );
  NAND2X1 U1607 ( .A(arr[783]), .B(n2747), .Y(n5320) );
  OAI21X1 U1608 ( .A(n4517), .B(n2746), .C(n5321), .Y(n7542) );
  NAND2X1 U1609 ( .A(arr[784]), .B(n2747), .Y(n5321) );
  OAI21X1 U1610 ( .A(n4519), .B(n2745), .C(n5322), .Y(n7543) );
  NAND2X1 U1611 ( .A(arr[785]), .B(n2746), .Y(n5322) );
  OAI21X1 U1612 ( .A(n4521), .B(n2746), .C(n5323), .Y(n7544) );
  NAND2X1 U1613 ( .A(arr[786]), .B(n2747), .Y(n5323) );
  OAI21X1 U1614 ( .A(n4523), .B(n2745), .C(n5324), .Y(n7545) );
  NAND2X1 U1615 ( .A(arr[787]), .B(n2746), .Y(n5324) );
  OAI21X1 U1616 ( .A(n4525), .B(n2745), .C(n5325), .Y(n7546) );
  NAND2X1 U1617 ( .A(arr[788]), .B(n2747), .Y(n5325) );
  OAI21X1 U1618 ( .A(n4527), .B(n2745), .C(n5326), .Y(n7547) );
  NAND2X1 U1619 ( .A(arr[789]), .B(n2746), .Y(n5326) );
  OAI21X1 U1620 ( .A(n4529), .B(n2745), .C(n5327), .Y(n7548) );
  NAND2X1 U1621 ( .A(arr[790]), .B(n2746), .Y(n5327) );
  OAI21X1 U1622 ( .A(n4531), .B(n2745), .C(n5328), .Y(n7549) );
  NAND2X1 U1623 ( .A(arr[791]), .B(n2747), .Y(n5328) );
  OAI21X1 U1625 ( .A(n4467), .B(n2742), .C(n5330), .Y(n7550) );
  NAND2X1 U1626 ( .A(arr[792]), .B(n2744), .Y(n5330) );
  OAI21X1 U1627 ( .A(n4469), .B(n2742), .C(n5331), .Y(n7551) );
  NAND2X1 U1628 ( .A(arr[793]), .B(n2744), .Y(n5331) );
  OAI21X1 U1629 ( .A(n4471), .B(n2742), .C(n5332), .Y(n7552) );
  NAND2X1 U1630 ( .A(arr[794]), .B(n2744), .Y(n5332) );
  OAI21X1 U1631 ( .A(n4473), .B(n2742), .C(n5333), .Y(n7553) );
  NAND2X1 U1632 ( .A(arr[795]), .B(n2744), .Y(n5333) );
  OAI21X1 U1633 ( .A(n4475), .B(n2743), .C(n5334), .Y(n7554) );
  NAND2X1 U1634 ( .A(arr[796]), .B(n2744), .Y(n5334) );
  OAI21X1 U1635 ( .A(n4477), .B(n2743), .C(n5335), .Y(n7555) );
  NAND2X1 U1636 ( .A(arr[797]), .B(n2743), .Y(n5335) );
  OAI21X1 U1637 ( .A(n4479), .B(n2743), .C(n5336), .Y(n7556) );
  NAND2X1 U1638 ( .A(arr[798]), .B(n2744), .Y(n5336) );
  OAI21X1 U1639 ( .A(n4481), .B(n2744), .C(n5337), .Y(n7557) );
  NAND2X1 U1640 ( .A(arr[799]), .B(n2744), .Y(n5337) );
  OAI21X1 U1641 ( .A(n4483), .B(n2743), .C(n5338), .Y(n7558) );
  NAND2X1 U1642 ( .A(arr[800]), .B(n2744), .Y(n5338) );
  OAI21X1 U1643 ( .A(n4485), .B(n2744), .C(n5339), .Y(n7559) );
  NAND2X1 U1644 ( .A(arr[801]), .B(n2742), .Y(n5339) );
  OAI21X1 U1645 ( .A(n4487), .B(n2744), .C(n5340), .Y(n7560) );
  NAND2X1 U1646 ( .A(arr[802]), .B(n2744), .Y(n5340) );
  OAI21X1 U1647 ( .A(n4489), .B(n2743), .C(n5341), .Y(n7561) );
  NAND2X1 U1648 ( .A(arr[803]), .B(n2742), .Y(n5341) );
  OAI21X1 U1649 ( .A(n4491), .B(n2744), .C(n5342), .Y(n7562) );
  NAND2X1 U1650 ( .A(arr[804]), .B(n2743), .Y(n5342) );
  OAI21X1 U1651 ( .A(n4493), .B(n2744), .C(n5343), .Y(n7563) );
  NAND2X1 U1652 ( .A(arr[805]), .B(n2743), .Y(n5343) );
  OAI21X1 U1653 ( .A(n4495), .B(n2743), .C(n5344), .Y(n7564) );
  NAND2X1 U1654 ( .A(arr[806]), .B(n2744), .Y(n5344) );
  OAI21X1 U1655 ( .A(n4497), .B(n2744), .C(n5345), .Y(n7565) );
  NAND2X1 U1656 ( .A(arr[807]), .B(n2742), .Y(n5345) );
  OAI21X1 U1657 ( .A(n4499), .B(n2744), .C(n5346), .Y(n7566) );
  NAND2X1 U1658 ( .A(arr[808]), .B(n2744), .Y(n5346) );
  OAI21X1 U1659 ( .A(n4501), .B(n2743), .C(n5347), .Y(n7567) );
  NAND2X1 U1660 ( .A(arr[809]), .B(n2742), .Y(n5347) );
  OAI21X1 U1661 ( .A(n4503), .B(n2743), .C(n5348), .Y(n7568) );
  NAND2X1 U1662 ( .A(arr[810]), .B(n2743), .Y(n5348) );
  OAI21X1 U1663 ( .A(n4505), .B(n2743), .C(n5349), .Y(n7569) );
  NAND2X1 U1664 ( .A(arr[811]), .B(n2744), .Y(n5349) );
  OAI21X1 U1665 ( .A(n4507), .B(n2743), .C(n5350), .Y(n7570) );
  NAND2X1 U1666 ( .A(arr[812]), .B(n2742), .Y(n5350) );
  OAI21X1 U1667 ( .A(n4509), .B(n2743), .C(n5351), .Y(n7571) );
  NAND2X1 U1668 ( .A(arr[813]), .B(n2743), .Y(n5351) );
  OAI21X1 U1669 ( .A(n4511), .B(n2743), .C(n5352), .Y(n7572) );
  NAND2X1 U1670 ( .A(arr[814]), .B(n2744), .Y(n5352) );
  OAI21X1 U1671 ( .A(n4513), .B(n2742), .C(n5353), .Y(n7573) );
  NAND2X1 U1672 ( .A(arr[815]), .B(n2744), .Y(n5353) );
  OAI21X1 U1673 ( .A(n4515), .B(n2743), .C(n5354), .Y(n7574) );
  NAND2X1 U1674 ( .A(arr[816]), .B(n2744), .Y(n5354) );
  OAI21X1 U1675 ( .A(n4517), .B(n2742), .C(n5355), .Y(n7575) );
  NAND2X1 U1676 ( .A(arr[817]), .B(n2743), .Y(n5355) );
  OAI21X1 U1677 ( .A(n4519), .B(n2742), .C(n5356), .Y(n7576) );
  NAND2X1 U1678 ( .A(arr[818]), .B(n2742), .Y(n5356) );
  OAI21X1 U1679 ( .A(n4521), .B(n2742), .C(n5357), .Y(n7577) );
  NAND2X1 U1680 ( .A(arr[819]), .B(n2744), .Y(n5357) );
  OAI21X1 U1681 ( .A(n4523), .B(n2742), .C(n5358), .Y(n7578) );
  NAND2X1 U1682 ( .A(arr[820]), .B(n2743), .Y(n5358) );
  OAI21X1 U1683 ( .A(n4525), .B(n2742), .C(n5359), .Y(n7579) );
  NAND2X1 U1684 ( .A(arr[821]), .B(n2743), .Y(n5359) );
  OAI21X1 U1685 ( .A(n4527), .B(n2742), .C(n5360), .Y(n7580) );
  NAND2X1 U1686 ( .A(arr[822]), .B(n2742), .Y(n5360) );
  OAI21X1 U1687 ( .A(n4529), .B(n2742), .C(n5361), .Y(n7581) );
  NAND2X1 U1688 ( .A(arr[823]), .B(n2744), .Y(n5361) );
  OAI21X1 U1689 ( .A(n4531), .B(n2742), .C(n5362), .Y(n7582) );
  NAND2X1 U1690 ( .A(arr[824]), .B(n2742), .Y(n5362) );
  OAI21X1 U1692 ( .A(n4467), .B(n2741), .C(n5365), .Y(n7583) );
  NAND2X1 U1693 ( .A(arr[825]), .B(n2740), .Y(n5365) );
  OAI21X1 U1694 ( .A(n4469), .B(n2739), .C(n5366), .Y(n7584) );
  NAND2X1 U1695 ( .A(arr[826]), .B(n2740), .Y(n5366) );
  OAI21X1 U1696 ( .A(n4471), .B(n2739), .C(n5367), .Y(n7585) );
  NAND2X1 U1697 ( .A(arr[827]), .B(n2740), .Y(n5367) );
  OAI21X1 U1698 ( .A(n4473), .B(n2739), .C(n5368), .Y(n7586) );
  NAND2X1 U1699 ( .A(arr[828]), .B(n2740), .Y(n5368) );
  OAI21X1 U1700 ( .A(n4475), .B(n2739), .C(n5369), .Y(n7587) );
  NAND2X1 U1701 ( .A(arr[829]), .B(n2740), .Y(n5369) );
  OAI21X1 U1702 ( .A(n4477), .B(n2739), .C(n5370), .Y(n7588) );
  NAND2X1 U1703 ( .A(arr[830]), .B(n2741), .Y(n5370) );
  OAI21X1 U1704 ( .A(n4479), .B(n2739), .C(n5371), .Y(n7589) );
  NAND2X1 U1705 ( .A(arr[831]), .B(n2741), .Y(n5371) );
  OAI21X1 U1706 ( .A(n4481), .B(n2740), .C(n5372), .Y(n7590) );
  NAND2X1 U1707 ( .A(arr[832]), .B(n2740), .Y(n5372) );
  OAI21X1 U1708 ( .A(n4483), .B(n2739), .C(n5373), .Y(n7591) );
  NAND2X1 U1709 ( .A(arr[833]), .B(n2740), .Y(n5373) );
  OAI21X1 U1710 ( .A(n4485), .B(n2740), .C(n5374), .Y(n7592) );
  NAND2X1 U1711 ( .A(arr[834]), .B(n2741), .Y(n5374) );
  OAI21X1 U1712 ( .A(n4487), .B(n2740), .C(n5375), .Y(n7593) );
  NAND2X1 U1713 ( .A(arr[835]), .B(n2741), .Y(n5375) );
  OAI21X1 U1714 ( .A(n4489), .B(n2739), .C(n5376), .Y(n7594) );
  NAND2X1 U1715 ( .A(arr[836]), .B(n2741), .Y(n5376) );
  OAI21X1 U1716 ( .A(n4491), .B(n2740), .C(n5377), .Y(n7595) );
  NAND2X1 U1717 ( .A(arr[837]), .B(n2741), .Y(n5377) );
  OAI21X1 U1718 ( .A(n4493), .B(n2740), .C(n5378), .Y(n7596) );
  NAND2X1 U1719 ( .A(arr[838]), .B(n2741), .Y(n5378) );
  OAI21X1 U1720 ( .A(n4495), .B(n2739), .C(n5379), .Y(n7597) );
  NAND2X1 U1721 ( .A(arr[839]), .B(n2741), .Y(n5379) );
  OAI21X1 U1722 ( .A(n4497), .B(n2740), .C(n5380), .Y(n7598) );
  NAND2X1 U1723 ( .A(arr[840]), .B(n2741), .Y(n5380) );
  OAI21X1 U1724 ( .A(n4499), .B(n2740), .C(n5381), .Y(n7599) );
  NAND2X1 U1725 ( .A(arr[841]), .B(n2741), .Y(n5381) );
  OAI21X1 U1726 ( .A(n4501), .B(n2739), .C(n5382), .Y(n7600) );
  NAND2X1 U1727 ( .A(arr[842]), .B(n2741), .Y(n5382) );
  OAI21X1 U1728 ( .A(n4503), .B(n2739), .C(n5383), .Y(n7601) );
  NAND2X1 U1729 ( .A(arr[843]), .B(n2741), .Y(n5383) );
  OAI21X1 U1730 ( .A(n4505), .B(n2739), .C(n5384), .Y(n7602) );
  NAND2X1 U1731 ( .A(arr[844]), .B(n2741), .Y(n5384) );
  OAI21X1 U1732 ( .A(n4507), .B(n2739), .C(n5385), .Y(n7603) );
  NAND2X1 U1733 ( .A(arr[845]), .B(n2741), .Y(n5385) );
  OAI21X1 U1734 ( .A(n4509), .B(n2739), .C(n5386), .Y(n7604) );
  NAND2X1 U1735 ( .A(arr[846]), .B(n2741), .Y(n5386) );
  OAI21X1 U1736 ( .A(n4511), .B(n2739), .C(n5387), .Y(n7605) );
  NAND2X1 U1737 ( .A(arr[847]), .B(n2741), .Y(n5387) );
  OAI21X1 U1738 ( .A(n4513), .B(n2741), .C(n5388), .Y(n7606) );
  NAND2X1 U1739 ( .A(arr[848]), .B(n2741), .Y(n5388) );
  OAI21X1 U1740 ( .A(n4515), .B(n2739), .C(n5389), .Y(n7607) );
  NAND2X1 U1741 ( .A(arr[849]), .B(n2741), .Y(n5389) );
  OAI21X1 U1742 ( .A(n4517), .B(n2740), .C(n5390), .Y(n7608) );
  NAND2X1 U1743 ( .A(arr[850]), .B(n2741), .Y(n5390) );
  OAI21X1 U1744 ( .A(n4519), .B(n2739), .C(n5391), .Y(n7609) );
  NAND2X1 U1745 ( .A(arr[851]), .B(n2740), .Y(n5391) );
  OAI21X1 U1746 ( .A(n4521), .B(n2740), .C(n5392), .Y(n7610) );
  NAND2X1 U1747 ( .A(arr[852]), .B(n2741), .Y(n5392) );
  OAI21X1 U1748 ( .A(n4523), .B(n2739), .C(n5393), .Y(n7611) );
  NAND2X1 U1749 ( .A(arr[853]), .B(n2740), .Y(n5393) );
  OAI21X1 U1750 ( .A(n4525), .B(n2739), .C(n5394), .Y(n7612) );
  NAND2X1 U1751 ( .A(arr[854]), .B(n2741), .Y(n5394) );
  OAI21X1 U1752 ( .A(n4527), .B(n2739), .C(n5395), .Y(n7613) );
  NAND2X1 U1753 ( .A(arr[855]), .B(n2740), .Y(n5395) );
  OAI21X1 U1754 ( .A(n4529), .B(n2739), .C(n5396), .Y(n7614) );
  NAND2X1 U1755 ( .A(arr[856]), .B(n2740), .Y(n5396) );
  OAI21X1 U1756 ( .A(n4531), .B(n2739), .C(n5397), .Y(n7615) );
  NAND2X1 U1757 ( .A(arr[857]), .B(n2741), .Y(n5397) );
  OAI21X1 U1759 ( .A(n4467), .B(n2736), .C(n5399), .Y(n7616) );
  NAND2X1 U1760 ( .A(arr[858]), .B(n2738), .Y(n5399) );
  OAI21X1 U1761 ( .A(n4469), .B(n2736), .C(n5400), .Y(n7617) );
  NAND2X1 U1762 ( .A(arr[859]), .B(n2738), .Y(n5400) );
  OAI21X1 U1763 ( .A(n4471), .B(n2736), .C(n5401), .Y(n7618) );
  NAND2X1 U1764 ( .A(arr[860]), .B(n2738), .Y(n5401) );
  OAI21X1 U1765 ( .A(n4473), .B(n2736), .C(n5402), .Y(n7619) );
  NAND2X1 U1766 ( .A(arr[861]), .B(n2738), .Y(n5402) );
  OAI21X1 U1767 ( .A(n4475), .B(n2737), .C(n5403), .Y(n7620) );
  NAND2X1 U1768 ( .A(arr[862]), .B(n2738), .Y(n5403) );
  OAI21X1 U1769 ( .A(n4477), .B(n2737), .C(n5404), .Y(n7621) );
  NAND2X1 U1770 ( .A(arr[863]), .B(n2737), .Y(n5404) );
  OAI21X1 U1771 ( .A(n4479), .B(n2737), .C(n5405), .Y(n7622) );
  NAND2X1 U1772 ( .A(arr[864]), .B(n2738), .Y(n5405) );
  OAI21X1 U1773 ( .A(n4481), .B(n2738), .C(n5406), .Y(n7623) );
  NAND2X1 U1774 ( .A(arr[865]), .B(n2738), .Y(n5406) );
  OAI21X1 U1775 ( .A(n4483), .B(n2737), .C(n5407), .Y(n7624) );
  NAND2X1 U1776 ( .A(arr[866]), .B(n2738), .Y(n5407) );
  OAI21X1 U1777 ( .A(n4485), .B(n2738), .C(n5408), .Y(n7625) );
  NAND2X1 U1778 ( .A(arr[867]), .B(n2736), .Y(n5408) );
  OAI21X1 U1779 ( .A(n4487), .B(n2738), .C(n5409), .Y(n7626) );
  NAND2X1 U1780 ( .A(arr[868]), .B(n2738), .Y(n5409) );
  OAI21X1 U1781 ( .A(n4489), .B(n2737), .C(n5410), .Y(n7627) );
  NAND2X1 U1782 ( .A(arr[869]), .B(n2736), .Y(n5410) );
  OAI21X1 U1783 ( .A(n4491), .B(n2738), .C(n5411), .Y(n7628) );
  NAND2X1 U1784 ( .A(arr[870]), .B(n2737), .Y(n5411) );
  OAI21X1 U1785 ( .A(n4493), .B(n2738), .C(n5412), .Y(n7629) );
  NAND2X1 U1786 ( .A(arr[871]), .B(n2737), .Y(n5412) );
  OAI21X1 U1787 ( .A(n4495), .B(n2737), .C(n5413), .Y(n7630) );
  NAND2X1 U1788 ( .A(arr[872]), .B(n2738), .Y(n5413) );
  OAI21X1 U1789 ( .A(n4497), .B(n2738), .C(n5414), .Y(n7631) );
  NAND2X1 U1790 ( .A(arr[873]), .B(n2736), .Y(n5414) );
  OAI21X1 U1791 ( .A(n4499), .B(n2738), .C(n5415), .Y(n7632) );
  NAND2X1 U1792 ( .A(arr[874]), .B(n2738), .Y(n5415) );
  OAI21X1 U1793 ( .A(n4501), .B(n2737), .C(n5416), .Y(n7633) );
  NAND2X1 U1794 ( .A(arr[875]), .B(n2736), .Y(n5416) );
  OAI21X1 U1795 ( .A(n4503), .B(n2737), .C(n5417), .Y(n7634) );
  NAND2X1 U1796 ( .A(arr[876]), .B(n2737), .Y(n5417) );
  OAI21X1 U1797 ( .A(n4505), .B(n2737), .C(n5418), .Y(n7635) );
  NAND2X1 U1798 ( .A(arr[877]), .B(n2738), .Y(n5418) );
  OAI21X1 U1799 ( .A(n4507), .B(n2737), .C(n5419), .Y(n7636) );
  NAND2X1 U1800 ( .A(arr[878]), .B(n2736), .Y(n5419) );
  OAI21X1 U1801 ( .A(n4509), .B(n2737), .C(n5420), .Y(n7637) );
  NAND2X1 U1802 ( .A(arr[879]), .B(n2737), .Y(n5420) );
  OAI21X1 U1803 ( .A(n4511), .B(n2737), .C(n5421), .Y(n7638) );
  NAND2X1 U1804 ( .A(arr[880]), .B(n2738), .Y(n5421) );
  OAI21X1 U1805 ( .A(n4513), .B(n2736), .C(n5422), .Y(n7639) );
  NAND2X1 U1806 ( .A(arr[881]), .B(n2738), .Y(n5422) );
  OAI21X1 U1807 ( .A(n4515), .B(n2737), .C(n5423), .Y(n7640) );
  NAND2X1 U1808 ( .A(arr[882]), .B(n2738), .Y(n5423) );
  OAI21X1 U1809 ( .A(n4517), .B(n2736), .C(n5424), .Y(n7641) );
  NAND2X1 U1810 ( .A(arr[883]), .B(n2737), .Y(n5424) );
  OAI21X1 U1811 ( .A(n4519), .B(n2736), .C(n5425), .Y(n7642) );
  NAND2X1 U1812 ( .A(arr[884]), .B(n2736), .Y(n5425) );
  OAI21X1 U1813 ( .A(n4521), .B(n2736), .C(n5426), .Y(n7643) );
  NAND2X1 U1814 ( .A(arr[885]), .B(n2738), .Y(n5426) );
  OAI21X1 U1815 ( .A(n4523), .B(n2736), .C(n5427), .Y(n7644) );
  NAND2X1 U1816 ( .A(arr[886]), .B(n2737), .Y(n5427) );
  OAI21X1 U1817 ( .A(n4525), .B(n2736), .C(n5428), .Y(n7645) );
  NAND2X1 U1818 ( .A(arr[887]), .B(n2737), .Y(n5428) );
  OAI21X1 U1819 ( .A(n4527), .B(n2736), .C(n5429), .Y(n7646) );
  NAND2X1 U1820 ( .A(arr[888]), .B(n2736), .Y(n5429) );
  OAI21X1 U1821 ( .A(n4529), .B(n2736), .C(n5430), .Y(n7647) );
  NAND2X1 U1822 ( .A(arr[889]), .B(n2738), .Y(n5430) );
  OAI21X1 U1823 ( .A(n4531), .B(n2736), .C(n5431), .Y(n7648) );
  NAND2X1 U1824 ( .A(arr[890]), .B(n2736), .Y(n5431) );
  OAI21X1 U1826 ( .A(n4467), .B(n2735), .C(n5434), .Y(n7649) );
  NAND2X1 U1827 ( .A(arr[891]), .B(n2734), .Y(n5434) );
  OAI21X1 U1828 ( .A(n4469), .B(n2733), .C(n5435), .Y(n7650) );
  NAND2X1 U1829 ( .A(arr[892]), .B(n2734), .Y(n5435) );
  OAI21X1 U1830 ( .A(n4471), .B(n2733), .C(n5436), .Y(n7651) );
  NAND2X1 U1831 ( .A(arr[893]), .B(n2734), .Y(n5436) );
  OAI21X1 U1832 ( .A(n4473), .B(n2733), .C(n5437), .Y(n7652) );
  NAND2X1 U1833 ( .A(arr[894]), .B(n2734), .Y(n5437) );
  OAI21X1 U1834 ( .A(n4475), .B(n2733), .C(n5438), .Y(n7653) );
  NAND2X1 U1835 ( .A(arr[895]), .B(n2734), .Y(n5438) );
  OAI21X1 U1836 ( .A(n4477), .B(n2733), .C(n5439), .Y(n7654) );
  NAND2X1 U1837 ( .A(arr[896]), .B(n2735), .Y(n5439) );
  OAI21X1 U1838 ( .A(n4479), .B(n2733), .C(n5440), .Y(n7655) );
  NAND2X1 U1839 ( .A(arr[897]), .B(n2735), .Y(n5440) );
  OAI21X1 U1840 ( .A(n4481), .B(n2734), .C(n5441), .Y(n7656) );
  NAND2X1 U1841 ( .A(arr[898]), .B(n2734), .Y(n5441) );
  OAI21X1 U1842 ( .A(n4483), .B(n2733), .C(n5442), .Y(n7657) );
  NAND2X1 U1843 ( .A(arr[899]), .B(n2734), .Y(n5442) );
  OAI21X1 U1844 ( .A(n4485), .B(n2734), .C(n5443), .Y(n7658) );
  NAND2X1 U1845 ( .A(arr[900]), .B(n2735), .Y(n5443) );
  OAI21X1 U1846 ( .A(n4487), .B(n2734), .C(n5444), .Y(n7659) );
  NAND2X1 U1847 ( .A(arr[901]), .B(n2735), .Y(n5444) );
  OAI21X1 U1848 ( .A(n4489), .B(n2733), .C(n5445), .Y(n7660) );
  NAND2X1 U1849 ( .A(arr[902]), .B(n2735), .Y(n5445) );
  OAI21X1 U1850 ( .A(n4491), .B(n2734), .C(n5446), .Y(n7661) );
  NAND2X1 U1851 ( .A(arr[903]), .B(n2735), .Y(n5446) );
  OAI21X1 U1852 ( .A(n4493), .B(n2734), .C(n5447), .Y(n7662) );
  NAND2X1 U1853 ( .A(arr[904]), .B(n2735), .Y(n5447) );
  OAI21X1 U1854 ( .A(n4495), .B(n2733), .C(n5448), .Y(n7663) );
  NAND2X1 U1855 ( .A(arr[905]), .B(n2735), .Y(n5448) );
  OAI21X1 U1856 ( .A(n4497), .B(n2734), .C(n5449), .Y(n7664) );
  NAND2X1 U1857 ( .A(arr[906]), .B(n2735), .Y(n5449) );
  OAI21X1 U1858 ( .A(n4499), .B(n2734), .C(n5450), .Y(n7665) );
  NAND2X1 U1859 ( .A(arr[907]), .B(n2735), .Y(n5450) );
  OAI21X1 U1860 ( .A(n4501), .B(n2733), .C(n5451), .Y(n7666) );
  NAND2X1 U1861 ( .A(arr[908]), .B(n2735), .Y(n5451) );
  OAI21X1 U1862 ( .A(n4503), .B(n2733), .C(n5452), .Y(n7667) );
  NAND2X1 U1863 ( .A(arr[909]), .B(n2735), .Y(n5452) );
  OAI21X1 U1864 ( .A(n4505), .B(n2733), .C(n5453), .Y(n7668) );
  NAND2X1 U1865 ( .A(arr[910]), .B(n2735), .Y(n5453) );
  OAI21X1 U1866 ( .A(n4507), .B(n2733), .C(n5454), .Y(n7669) );
  NAND2X1 U1867 ( .A(arr[911]), .B(n2735), .Y(n5454) );
  OAI21X1 U1868 ( .A(n4509), .B(n2733), .C(n5455), .Y(n7670) );
  NAND2X1 U1869 ( .A(arr[912]), .B(n2735), .Y(n5455) );
  OAI21X1 U1870 ( .A(n4511), .B(n2733), .C(n5456), .Y(n7671) );
  NAND2X1 U1871 ( .A(arr[913]), .B(n2735), .Y(n5456) );
  OAI21X1 U1872 ( .A(n4513), .B(n2735), .C(n5457), .Y(n7672) );
  NAND2X1 U1873 ( .A(arr[914]), .B(n2735), .Y(n5457) );
  OAI21X1 U1874 ( .A(n4515), .B(n2733), .C(n5458), .Y(n7673) );
  NAND2X1 U1875 ( .A(arr[915]), .B(n2735), .Y(n5458) );
  OAI21X1 U1876 ( .A(n4517), .B(n2734), .C(n5459), .Y(n7674) );
  NAND2X1 U1877 ( .A(arr[916]), .B(n2735), .Y(n5459) );
  OAI21X1 U1878 ( .A(n4519), .B(n2733), .C(n5460), .Y(n7675) );
  NAND2X1 U1879 ( .A(arr[917]), .B(n2734), .Y(n5460) );
  OAI21X1 U1880 ( .A(n4521), .B(n2734), .C(n5461), .Y(n7676) );
  NAND2X1 U1881 ( .A(arr[918]), .B(n2735), .Y(n5461) );
  OAI21X1 U1882 ( .A(n4523), .B(n2733), .C(n5462), .Y(n7677) );
  NAND2X1 U1883 ( .A(arr[919]), .B(n2734), .Y(n5462) );
  OAI21X1 U1884 ( .A(n4525), .B(n2733), .C(n5463), .Y(n7678) );
  NAND2X1 U1885 ( .A(arr[920]), .B(n2735), .Y(n5463) );
  OAI21X1 U1886 ( .A(n4527), .B(n2733), .C(n5464), .Y(n7679) );
  NAND2X1 U1887 ( .A(arr[921]), .B(n2734), .Y(n5464) );
  OAI21X1 U1888 ( .A(n4529), .B(n2733), .C(n5465), .Y(n7680) );
  NAND2X1 U1889 ( .A(arr[922]), .B(n2734), .Y(n5465) );
  OAI21X1 U1890 ( .A(n4531), .B(n2733), .C(n5466), .Y(n7681) );
  NAND2X1 U1891 ( .A(arr[923]), .B(n2735), .Y(n5466) );
  OAI21X1 U1893 ( .A(n4467), .B(n2730), .C(n5468), .Y(n7682) );
  NAND2X1 U1894 ( .A(arr[924]), .B(n2732), .Y(n5468) );
  OAI21X1 U1895 ( .A(n4469), .B(n2730), .C(n5469), .Y(n7683) );
  NAND2X1 U1896 ( .A(arr[925]), .B(n2732), .Y(n5469) );
  OAI21X1 U1897 ( .A(n4471), .B(n2730), .C(n5470), .Y(n7684) );
  NAND2X1 U1898 ( .A(arr[926]), .B(n2732), .Y(n5470) );
  OAI21X1 U1899 ( .A(n4473), .B(n2730), .C(n5471), .Y(n7685) );
  NAND2X1 U1900 ( .A(arr[927]), .B(n2732), .Y(n5471) );
  OAI21X1 U1901 ( .A(n4475), .B(n2731), .C(n5472), .Y(n7686) );
  NAND2X1 U1902 ( .A(arr[928]), .B(n2732), .Y(n5472) );
  OAI21X1 U1903 ( .A(n4477), .B(n2731), .C(n5473), .Y(n7687) );
  NAND2X1 U1904 ( .A(arr[929]), .B(n2731), .Y(n5473) );
  OAI21X1 U1905 ( .A(n4479), .B(n2731), .C(n5474), .Y(n7688) );
  NAND2X1 U1906 ( .A(arr[930]), .B(n2732), .Y(n5474) );
  OAI21X1 U1907 ( .A(n4481), .B(n2732), .C(n5475), .Y(n7689) );
  NAND2X1 U1908 ( .A(arr[931]), .B(n2732), .Y(n5475) );
  OAI21X1 U1909 ( .A(n4483), .B(n2731), .C(n5476), .Y(n7690) );
  NAND2X1 U1910 ( .A(arr[932]), .B(n2732), .Y(n5476) );
  OAI21X1 U1911 ( .A(n4485), .B(n2732), .C(n5477), .Y(n7691) );
  NAND2X1 U1912 ( .A(arr[933]), .B(n2730), .Y(n5477) );
  OAI21X1 U1913 ( .A(n4487), .B(n2732), .C(n5478), .Y(n7692) );
  NAND2X1 U1914 ( .A(arr[934]), .B(n2732), .Y(n5478) );
  OAI21X1 U1915 ( .A(n4489), .B(n2731), .C(n5479), .Y(n7693) );
  NAND2X1 U1916 ( .A(arr[935]), .B(n2730), .Y(n5479) );
  OAI21X1 U1917 ( .A(n4491), .B(n2732), .C(n5480), .Y(n7694) );
  NAND2X1 U1918 ( .A(arr[936]), .B(n2731), .Y(n5480) );
  OAI21X1 U1919 ( .A(n4493), .B(n2732), .C(n5481), .Y(n7695) );
  NAND2X1 U1920 ( .A(arr[937]), .B(n2731), .Y(n5481) );
  OAI21X1 U1921 ( .A(n4495), .B(n2731), .C(n5482), .Y(n7696) );
  NAND2X1 U1922 ( .A(arr[938]), .B(n2732), .Y(n5482) );
  OAI21X1 U1923 ( .A(n4497), .B(n2732), .C(n5483), .Y(n7697) );
  NAND2X1 U1924 ( .A(arr[939]), .B(n2730), .Y(n5483) );
  OAI21X1 U1925 ( .A(n4499), .B(n2732), .C(n5484), .Y(n7698) );
  NAND2X1 U1926 ( .A(arr[940]), .B(n2732), .Y(n5484) );
  OAI21X1 U1927 ( .A(n4501), .B(n2731), .C(n5485), .Y(n7699) );
  NAND2X1 U1928 ( .A(arr[941]), .B(n2730), .Y(n5485) );
  OAI21X1 U1929 ( .A(n4503), .B(n2731), .C(n5486), .Y(n7700) );
  NAND2X1 U1930 ( .A(arr[942]), .B(n2731), .Y(n5486) );
  OAI21X1 U1931 ( .A(n4505), .B(n2731), .C(n5487), .Y(n7701) );
  NAND2X1 U1932 ( .A(arr[943]), .B(n2732), .Y(n5487) );
  OAI21X1 U1933 ( .A(n4507), .B(n2731), .C(n5488), .Y(n7702) );
  NAND2X1 U1934 ( .A(arr[944]), .B(n2730), .Y(n5488) );
  OAI21X1 U1935 ( .A(n4509), .B(n2731), .C(n5489), .Y(n7703) );
  NAND2X1 U1936 ( .A(arr[945]), .B(n2731), .Y(n5489) );
  OAI21X1 U1937 ( .A(n4511), .B(n2731), .C(n5490), .Y(n7704) );
  NAND2X1 U1938 ( .A(arr[946]), .B(n2732), .Y(n5490) );
  OAI21X1 U1939 ( .A(n4513), .B(n2730), .C(n5491), .Y(n7705) );
  NAND2X1 U1940 ( .A(arr[947]), .B(n2732), .Y(n5491) );
  OAI21X1 U1941 ( .A(n4515), .B(n2731), .C(n5492), .Y(n7706) );
  NAND2X1 U1942 ( .A(arr[948]), .B(n2732), .Y(n5492) );
  OAI21X1 U1943 ( .A(n4517), .B(n2730), .C(n5493), .Y(n7707) );
  NAND2X1 U1944 ( .A(arr[949]), .B(n2731), .Y(n5493) );
  OAI21X1 U1945 ( .A(n4519), .B(n2730), .C(n5494), .Y(n7708) );
  NAND2X1 U1946 ( .A(arr[950]), .B(n2730), .Y(n5494) );
  OAI21X1 U1947 ( .A(n4521), .B(n2730), .C(n5495), .Y(n7709) );
  NAND2X1 U1948 ( .A(arr[951]), .B(n2732), .Y(n5495) );
  OAI21X1 U1949 ( .A(n4523), .B(n2730), .C(n5496), .Y(n7710) );
  NAND2X1 U1950 ( .A(arr[952]), .B(n2731), .Y(n5496) );
  OAI21X1 U1951 ( .A(n4525), .B(n2730), .C(n5497), .Y(n7711) );
  NAND2X1 U1952 ( .A(arr[953]), .B(n2731), .Y(n5497) );
  OAI21X1 U1953 ( .A(n4527), .B(n2730), .C(n5498), .Y(n7712) );
  NAND2X1 U1954 ( .A(arr[954]), .B(n2730), .Y(n5498) );
  OAI21X1 U1955 ( .A(n4529), .B(n2730), .C(n5499), .Y(n7713) );
  NAND2X1 U1956 ( .A(arr[955]), .B(n2732), .Y(n5499) );
  OAI21X1 U1957 ( .A(n4531), .B(n2730), .C(n5500), .Y(n7714) );
  NAND2X1 U1958 ( .A(arr[956]), .B(n2730), .Y(n5500) );
  OAI21X1 U1960 ( .A(n4467), .B(n2729), .C(n5503), .Y(n7715) );
  NAND2X1 U1961 ( .A(arr[957]), .B(n2728), .Y(n5503) );
  OAI21X1 U1962 ( .A(n4469), .B(n2727), .C(n5504), .Y(n7716) );
  NAND2X1 U1963 ( .A(arr[958]), .B(n2728), .Y(n5504) );
  OAI21X1 U1964 ( .A(n4471), .B(n2727), .C(n5505), .Y(n7717) );
  NAND2X1 U1965 ( .A(arr[959]), .B(n2728), .Y(n5505) );
  OAI21X1 U1966 ( .A(n4473), .B(n2727), .C(n5506), .Y(n7718) );
  NAND2X1 U1967 ( .A(arr[960]), .B(n2728), .Y(n5506) );
  OAI21X1 U1968 ( .A(n4475), .B(n2727), .C(n5507), .Y(n7719) );
  NAND2X1 U1969 ( .A(arr[961]), .B(n2728), .Y(n5507) );
  OAI21X1 U1970 ( .A(n4477), .B(n2727), .C(n5508), .Y(n7720) );
  NAND2X1 U1971 ( .A(arr[962]), .B(n2729), .Y(n5508) );
  OAI21X1 U1972 ( .A(n4479), .B(n2727), .C(n5509), .Y(n7721) );
  NAND2X1 U1973 ( .A(arr[963]), .B(n2729), .Y(n5509) );
  OAI21X1 U1974 ( .A(n4481), .B(n2728), .C(n5510), .Y(n7722) );
  NAND2X1 U1975 ( .A(arr[964]), .B(n2728), .Y(n5510) );
  OAI21X1 U1976 ( .A(n4483), .B(n2727), .C(n5511), .Y(n7723) );
  NAND2X1 U1977 ( .A(arr[965]), .B(n2728), .Y(n5511) );
  OAI21X1 U1978 ( .A(n4485), .B(n2728), .C(n5512), .Y(n7724) );
  NAND2X1 U1979 ( .A(arr[966]), .B(n2729), .Y(n5512) );
  OAI21X1 U1980 ( .A(n4487), .B(n2728), .C(n5513), .Y(n7725) );
  NAND2X1 U1981 ( .A(arr[967]), .B(n2729), .Y(n5513) );
  OAI21X1 U1982 ( .A(n4489), .B(n2727), .C(n5514), .Y(n7726) );
  NAND2X1 U1983 ( .A(arr[968]), .B(n2729), .Y(n5514) );
  OAI21X1 U1984 ( .A(n4491), .B(n2728), .C(n5515), .Y(n7727) );
  NAND2X1 U1985 ( .A(arr[969]), .B(n2729), .Y(n5515) );
  OAI21X1 U1986 ( .A(n4493), .B(n2728), .C(n5516), .Y(n7728) );
  NAND2X1 U1987 ( .A(arr[970]), .B(n2729), .Y(n5516) );
  OAI21X1 U1988 ( .A(n4495), .B(n2727), .C(n5517), .Y(n7729) );
  NAND2X1 U1989 ( .A(arr[971]), .B(n2729), .Y(n5517) );
  OAI21X1 U1990 ( .A(n4497), .B(n2728), .C(n5518), .Y(n7730) );
  NAND2X1 U1991 ( .A(arr[972]), .B(n2729), .Y(n5518) );
  OAI21X1 U1992 ( .A(n4499), .B(n2728), .C(n5519), .Y(n7731) );
  NAND2X1 U1993 ( .A(arr[973]), .B(n2729), .Y(n5519) );
  OAI21X1 U1994 ( .A(n4501), .B(n2727), .C(n5520), .Y(n7732) );
  NAND2X1 U1995 ( .A(arr[974]), .B(n2729), .Y(n5520) );
  OAI21X1 U1996 ( .A(n4503), .B(n2727), .C(n5521), .Y(n7733) );
  NAND2X1 U1997 ( .A(arr[975]), .B(n2729), .Y(n5521) );
  OAI21X1 U1998 ( .A(n4505), .B(n2727), .C(n5522), .Y(n7734) );
  NAND2X1 U1999 ( .A(arr[976]), .B(n2729), .Y(n5522) );
  OAI21X1 U2000 ( .A(n4507), .B(n2727), .C(n5523), .Y(n7735) );
  NAND2X1 U2001 ( .A(arr[977]), .B(n2729), .Y(n5523) );
  OAI21X1 U2002 ( .A(n4509), .B(n2727), .C(n5524), .Y(n7736) );
  NAND2X1 U2003 ( .A(arr[978]), .B(n2729), .Y(n5524) );
  OAI21X1 U2004 ( .A(n4511), .B(n2727), .C(n5525), .Y(n7737) );
  NAND2X1 U2005 ( .A(arr[979]), .B(n2729), .Y(n5525) );
  OAI21X1 U2006 ( .A(n4513), .B(n2729), .C(n5526), .Y(n7738) );
  NAND2X1 U2007 ( .A(arr[980]), .B(n2729), .Y(n5526) );
  OAI21X1 U2008 ( .A(n4515), .B(n2727), .C(n5527), .Y(n7739) );
  NAND2X1 U2009 ( .A(arr[981]), .B(n2729), .Y(n5527) );
  OAI21X1 U2010 ( .A(n4517), .B(n2728), .C(n5528), .Y(n7740) );
  NAND2X1 U2011 ( .A(arr[982]), .B(n2729), .Y(n5528) );
  OAI21X1 U2012 ( .A(n4519), .B(n2727), .C(n5529), .Y(n7741) );
  NAND2X1 U2013 ( .A(arr[983]), .B(n2728), .Y(n5529) );
  OAI21X1 U2014 ( .A(n4521), .B(n2728), .C(n5530), .Y(n7742) );
  NAND2X1 U2015 ( .A(arr[984]), .B(n2729), .Y(n5530) );
  OAI21X1 U2016 ( .A(n4523), .B(n2727), .C(n5531), .Y(n7743) );
  NAND2X1 U2017 ( .A(arr[985]), .B(n2728), .Y(n5531) );
  OAI21X1 U2018 ( .A(n4525), .B(n2727), .C(n5532), .Y(n7744) );
  NAND2X1 U2019 ( .A(arr[986]), .B(n2729), .Y(n5532) );
  OAI21X1 U2020 ( .A(n4527), .B(n2727), .C(n5533), .Y(n7745) );
  NAND2X1 U2021 ( .A(arr[987]), .B(n2728), .Y(n5533) );
  OAI21X1 U2022 ( .A(n4529), .B(n2727), .C(n5534), .Y(n7746) );
  NAND2X1 U2023 ( .A(arr[988]), .B(n2728), .Y(n5534) );
  OAI21X1 U2024 ( .A(n4531), .B(n2727), .C(n5535), .Y(n7747) );
  NAND2X1 U2025 ( .A(arr[989]), .B(n2729), .Y(n5535) );
  OAI21X1 U2027 ( .A(n4467), .B(n2724), .C(n5537), .Y(n7748) );
  NAND2X1 U2028 ( .A(arr[990]), .B(n2726), .Y(n5537) );
  OAI21X1 U2029 ( .A(n4469), .B(n2724), .C(n5538), .Y(n7749) );
  NAND2X1 U2030 ( .A(arr[991]), .B(n2726), .Y(n5538) );
  OAI21X1 U2031 ( .A(n4471), .B(n2724), .C(n5539), .Y(n7750) );
  NAND2X1 U2032 ( .A(arr[992]), .B(n2726), .Y(n5539) );
  OAI21X1 U2033 ( .A(n4473), .B(n2724), .C(n5540), .Y(n7751) );
  NAND2X1 U2034 ( .A(arr[993]), .B(n2726), .Y(n5540) );
  OAI21X1 U2035 ( .A(n4475), .B(n2725), .C(n5541), .Y(n7752) );
  NAND2X1 U2036 ( .A(arr[994]), .B(n2726), .Y(n5541) );
  OAI21X1 U2037 ( .A(n4477), .B(n2725), .C(n5542), .Y(n7753) );
  NAND2X1 U2038 ( .A(arr[995]), .B(n2725), .Y(n5542) );
  OAI21X1 U2039 ( .A(n4479), .B(n2725), .C(n5543), .Y(n7754) );
  NAND2X1 U2040 ( .A(arr[996]), .B(n2726), .Y(n5543) );
  OAI21X1 U2041 ( .A(n4481), .B(n2726), .C(n5544), .Y(n7755) );
  NAND2X1 U2042 ( .A(arr[997]), .B(n2726), .Y(n5544) );
  OAI21X1 U2043 ( .A(n4483), .B(n2725), .C(n5545), .Y(n7756) );
  NAND2X1 U2044 ( .A(arr[998]), .B(n2726), .Y(n5545) );
  OAI21X1 U2045 ( .A(n4485), .B(n2726), .C(n5546), .Y(n7757) );
  NAND2X1 U2046 ( .A(arr[999]), .B(n2724), .Y(n5546) );
  OAI21X1 U2047 ( .A(n4487), .B(n2726), .C(n5547), .Y(n7758) );
  NAND2X1 U2048 ( .A(arr[1000]), .B(n2726), .Y(n5547) );
  OAI21X1 U2049 ( .A(n4489), .B(n2725), .C(n5548), .Y(n7759) );
  NAND2X1 U2050 ( .A(arr[1001]), .B(n2724), .Y(n5548) );
  OAI21X1 U2051 ( .A(n4491), .B(n2726), .C(n5549), .Y(n7760) );
  NAND2X1 U2052 ( .A(arr[1002]), .B(n2725), .Y(n5549) );
  OAI21X1 U2053 ( .A(n4493), .B(n2726), .C(n5550), .Y(n7761) );
  NAND2X1 U2054 ( .A(arr[1003]), .B(n2725), .Y(n5550) );
  OAI21X1 U2055 ( .A(n4495), .B(n2725), .C(n5551), .Y(n7762) );
  NAND2X1 U2056 ( .A(arr[1004]), .B(n2726), .Y(n5551) );
  OAI21X1 U2057 ( .A(n4497), .B(n2726), .C(n5552), .Y(n7763) );
  NAND2X1 U2058 ( .A(arr[1005]), .B(n2724), .Y(n5552) );
  OAI21X1 U2059 ( .A(n4499), .B(n2726), .C(n5553), .Y(n7764) );
  NAND2X1 U2060 ( .A(arr[1006]), .B(n2726), .Y(n5553) );
  OAI21X1 U2061 ( .A(n4501), .B(n2725), .C(n5554), .Y(n7765) );
  NAND2X1 U2062 ( .A(arr[1007]), .B(n2724), .Y(n5554) );
  OAI21X1 U2063 ( .A(n4503), .B(n2725), .C(n5555), .Y(n7766) );
  NAND2X1 U2064 ( .A(arr[1008]), .B(n2725), .Y(n5555) );
  OAI21X1 U2065 ( .A(n4505), .B(n2725), .C(n5556), .Y(n7767) );
  NAND2X1 U2066 ( .A(arr[1009]), .B(n2726), .Y(n5556) );
  OAI21X1 U2067 ( .A(n4507), .B(n2725), .C(n5557), .Y(n7768) );
  NAND2X1 U2068 ( .A(arr[1010]), .B(n2724), .Y(n5557) );
  OAI21X1 U2069 ( .A(n4509), .B(n2725), .C(n5558), .Y(n7769) );
  NAND2X1 U2070 ( .A(arr[1011]), .B(n2725), .Y(n5558) );
  OAI21X1 U2071 ( .A(n4511), .B(n2725), .C(n5559), .Y(n7770) );
  NAND2X1 U2072 ( .A(arr[1012]), .B(n2726), .Y(n5559) );
  OAI21X1 U2073 ( .A(n4513), .B(n2724), .C(n5560), .Y(n7771) );
  NAND2X1 U2074 ( .A(arr[1013]), .B(n2726), .Y(n5560) );
  OAI21X1 U2075 ( .A(n4515), .B(n2725), .C(n5561), .Y(n7772) );
  NAND2X1 U2076 ( .A(arr[1014]), .B(n2726), .Y(n5561) );
  OAI21X1 U2077 ( .A(n4517), .B(n2724), .C(n5562), .Y(n7773) );
  NAND2X1 U2078 ( .A(arr[1015]), .B(n2725), .Y(n5562) );
  OAI21X1 U2079 ( .A(n4519), .B(n2724), .C(n5563), .Y(n7774) );
  NAND2X1 U2080 ( .A(arr[1016]), .B(n2724), .Y(n5563) );
  OAI21X1 U2081 ( .A(n4521), .B(n2724), .C(n5564), .Y(n7775) );
  NAND2X1 U2082 ( .A(arr[1017]), .B(n2726), .Y(n5564) );
  OAI21X1 U2083 ( .A(n4523), .B(n2724), .C(n5565), .Y(n7776) );
  NAND2X1 U2084 ( .A(arr[1018]), .B(n2725), .Y(n5565) );
  OAI21X1 U2085 ( .A(n4525), .B(n2724), .C(n5566), .Y(n7777) );
  NAND2X1 U2086 ( .A(arr[1019]), .B(n2725), .Y(n5566) );
  OAI21X1 U2087 ( .A(n4527), .B(n2724), .C(n5567), .Y(n7778) );
  NAND2X1 U2088 ( .A(arr[1020]), .B(n2724), .Y(n5567) );
  OAI21X1 U2089 ( .A(n4529), .B(n2724), .C(n5568), .Y(n7779) );
  NAND2X1 U2090 ( .A(arr[1021]), .B(n2726), .Y(n5568) );
  OAI21X1 U2091 ( .A(n4531), .B(n2724), .C(n5569), .Y(n7780) );
  NAND2X1 U2092 ( .A(arr[1022]), .B(n2724), .Y(n5569) );
  OAI21X1 U2095 ( .A(n4467), .B(n2723), .C(n5574), .Y(n7781) );
  NAND2X1 U2096 ( .A(arr[1023]), .B(n2722), .Y(n5574) );
  OAI21X1 U2097 ( .A(n4469), .B(n2721), .C(n5575), .Y(n7782) );
  NAND2X1 U2098 ( .A(arr[1024]), .B(n2722), .Y(n5575) );
  OAI21X1 U2099 ( .A(n4471), .B(n2721), .C(n5576), .Y(n7783) );
  NAND2X1 U2100 ( .A(arr[1025]), .B(n2722), .Y(n5576) );
  OAI21X1 U2101 ( .A(n4473), .B(n2721), .C(n5577), .Y(n7784) );
  NAND2X1 U2102 ( .A(arr[1026]), .B(n2722), .Y(n5577) );
  OAI21X1 U2103 ( .A(n4475), .B(n2721), .C(n5578), .Y(n7785) );
  NAND2X1 U2104 ( .A(arr[1027]), .B(n2722), .Y(n5578) );
  OAI21X1 U2105 ( .A(n4477), .B(n2721), .C(n5579), .Y(n7786) );
  NAND2X1 U2106 ( .A(arr[1028]), .B(n2723), .Y(n5579) );
  OAI21X1 U2107 ( .A(n4479), .B(n2721), .C(n5580), .Y(n7787) );
  NAND2X1 U2108 ( .A(arr[1029]), .B(n2723), .Y(n5580) );
  OAI21X1 U2109 ( .A(n4481), .B(n2722), .C(n5581), .Y(n7788) );
  NAND2X1 U2110 ( .A(arr[1030]), .B(n2722), .Y(n5581) );
  OAI21X1 U2111 ( .A(n4483), .B(n2721), .C(n5582), .Y(n7789) );
  NAND2X1 U2112 ( .A(arr[1031]), .B(n2722), .Y(n5582) );
  OAI21X1 U2113 ( .A(n4485), .B(n2722), .C(n5583), .Y(n7790) );
  NAND2X1 U2114 ( .A(arr[1032]), .B(n2723), .Y(n5583) );
  OAI21X1 U2115 ( .A(n4487), .B(n2722), .C(n5584), .Y(n7791) );
  NAND2X1 U2116 ( .A(arr[1033]), .B(n2723), .Y(n5584) );
  OAI21X1 U2117 ( .A(n4489), .B(n2721), .C(n5585), .Y(n7792) );
  NAND2X1 U2118 ( .A(arr[1034]), .B(n2723), .Y(n5585) );
  OAI21X1 U2119 ( .A(n4491), .B(n2722), .C(n5586), .Y(n7793) );
  NAND2X1 U2120 ( .A(arr[1035]), .B(n2723), .Y(n5586) );
  OAI21X1 U2121 ( .A(n4493), .B(n2722), .C(n5587), .Y(n7794) );
  NAND2X1 U2122 ( .A(arr[1036]), .B(n2723), .Y(n5587) );
  OAI21X1 U2123 ( .A(n4495), .B(n2721), .C(n5588), .Y(n7795) );
  NAND2X1 U2124 ( .A(arr[1037]), .B(n2723), .Y(n5588) );
  OAI21X1 U2125 ( .A(n4497), .B(n2722), .C(n5589), .Y(n7796) );
  NAND2X1 U2126 ( .A(arr[1038]), .B(n2723), .Y(n5589) );
  OAI21X1 U2127 ( .A(n4499), .B(n2722), .C(n5590), .Y(n7797) );
  NAND2X1 U2128 ( .A(arr[1039]), .B(n2723), .Y(n5590) );
  OAI21X1 U2129 ( .A(n4501), .B(n2721), .C(n5591), .Y(n7798) );
  NAND2X1 U2130 ( .A(arr[1040]), .B(n2723), .Y(n5591) );
  OAI21X1 U2131 ( .A(n4503), .B(n2721), .C(n5592), .Y(n7799) );
  NAND2X1 U2132 ( .A(arr[1041]), .B(n2723), .Y(n5592) );
  OAI21X1 U2133 ( .A(n4505), .B(n2721), .C(n5593), .Y(n7800) );
  NAND2X1 U2134 ( .A(arr[1042]), .B(n2723), .Y(n5593) );
  OAI21X1 U2135 ( .A(n4507), .B(n2721), .C(n5594), .Y(n7801) );
  NAND2X1 U2136 ( .A(arr[1043]), .B(n2723), .Y(n5594) );
  OAI21X1 U2137 ( .A(n4509), .B(n2721), .C(n5595), .Y(n7802) );
  NAND2X1 U2138 ( .A(arr[1044]), .B(n2723), .Y(n5595) );
  OAI21X1 U2139 ( .A(n4511), .B(n2721), .C(n5596), .Y(n7803) );
  NAND2X1 U2140 ( .A(arr[1045]), .B(n2723), .Y(n5596) );
  OAI21X1 U2141 ( .A(n4513), .B(n2723), .C(n5597), .Y(n7804) );
  NAND2X1 U2142 ( .A(arr[1046]), .B(n2723), .Y(n5597) );
  OAI21X1 U2143 ( .A(n4515), .B(n2721), .C(n5598), .Y(n7805) );
  NAND2X1 U2144 ( .A(arr[1047]), .B(n2723), .Y(n5598) );
  OAI21X1 U2145 ( .A(n4517), .B(n2722), .C(n5599), .Y(n7806) );
  NAND2X1 U2146 ( .A(arr[1048]), .B(n2723), .Y(n5599) );
  OAI21X1 U2147 ( .A(n4519), .B(n2721), .C(n5600), .Y(n7807) );
  NAND2X1 U2148 ( .A(arr[1049]), .B(n2722), .Y(n5600) );
  OAI21X1 U2149 ( .A(n4521), .B(n2722), .C(n5601), .Y(n7808) );
  NAND2X1 U2150 ( .A(arr[1050]), .B(n2723), .Y(n5601) );
  OAI21X1 U2151 ( .A(n4523), .B(n2721), .C(n5602), .Y(n7809) );
  NAND2X1 U2152 ( .A(arr[1051]), .B(n2722), .Y(n5602) );
  OAI21X1 U2153 ( .A(n4525), .B(n2721), .C(n5603), .Y(n7810) );
  NAND2X1 U2154 ( .A(arr[1052]), .B(n2723), .Y(n5603) );
  OAI21X1 U2155 ( .A(n4527), .B(n2721), .C(n5604), .Y(n7811) );
  NAND2X1 U2156 ( .A(arr[1053]), .B(n2722), .Y(n5604) );
  OAI21X1 U2157 ( .A(n4529), .B(n2721), .C(n5605), .Y(n7812) );
  NAND2X1 U2158 ( .A(arr[1054]), .B(n2722), .Y(n5605) );
  OAI21X1 U2159 ( .A(n4531), .B(n2721), .C(n5606), .Y(n7813) );
  NAND2X1 U2160 ( .A(arr[1055]), .B(n2723), .Y(n5606) );
  AND2X1 U2163 ( .A(n5607), .B(n5608), .Y(n5571) );
  OAI21X1 U2164 ( .A(n4467), .B(n2720), .C(n5610), .Y(n7814) );
  NAND2X1 U2165 ( .A(arr[1056]), .B(n2719), .Y(n5610) );
  OAI21X1 U2166 ( .A(n4469), .B(n2718), .C(n5611), .Y(n7815) );
  NAND2X1 U2167 ( .A(arr[1057]), .B(n2719), .Y(n5611) );
  OAI21X1 U2168 ( .A(n4471), .B(n2718), .C(n5612), .Y(n7816) );
  NAND2X1 U2169 ( .A(arr[1058]), .B(n2719), .Y(n5612) );
  OAI21X1 U2170 ( .A(n4473), .B(n2718), .C(n5613), .Y(n7817) );
  NAND2X1 U2171 ( .A(arr[1059]), .B(n2719), .Y(n5613) );
  OAI21X1 U2172 ( .A(n4475), .B(n2718), .C(n5614), .Y(n7818) );
  NAND2X1 U2173 ( .A(arr[1060]), .B(n2719), .Y(n5614) );
  OAI21X1 U2174 ( .A(n4477), .B(n2718), .C(n5615), .Y(n7819) );
  NAND2X1 U2175 ( .A(arr[1061]), .B(n2720), .Y(n5615) );
  OAI21X1 U2176 ( .A(n4479), .B(n2718), .C(n5616), .Y(n7820) );
  NAND2X1 U2177 ( .A(arr[1062]), .B(n2720), .Y(n5616) );
  OAI21X1 U2178 ( .A(n4481), .B(n2719), .C(n5617), .Y(n7821) );
  NAND2X1 U2179 ( .A(arr[1063]), .B(n2719), .Y(n5617) );
  OAI21X1 U2180 ( .A(n4483), .B(n2718), .C(n5618), .Y(n7822) );
  NAND2X1 U2181 ( .A(arr[1064]), .B(n2719), .Y(n5618) );
  OAI21X1 U2182 ( .A(n4485), .B(n2719), .C(n5619), .Y(n7823) );
  NAND2X1 U2183 ( .A(arr[1065]), .B(n2720), .Y(n5619) );
  OAI21X1 U2184 ( .A(n4487), .B(n2719), .C(n5620), .Y(n7824) );
  NAND2X1 U2185 ( .A(arr[1066]), .B(n2720), .Y(n5620) );
  OAI21X1 U2186 ( .A(n4489), .B(n2718), .C(n5621), .Y(n7825) );
  NAND2X1 U2187 ( .A(arr[1067]), .B(n2720), .Y(n5621) );
  OAI21X1 U2188 ( .A(n4491), .B(n2719), .C(n5622), .Y(n7826) );
  NAND2X1 U2189 ( .A(arr[1068]), .B(n2720), .Y(n5622) );
  OAI21X1 U2190 ( .A(n4493), .B(n2719), .C(n5623), .Y(n7827) );
  NAND2X1 U2191 ( .A(arr[1069]), .B(n2720), .Y(n5623) );
  OAI21X1 U2192 ( .A(n4495), .B(n2718), .C(n5624), .Y(n7828) );
  NAND2X1 U2193 ( .A(arr[1070]), .B(n2720), .Y(n5624) );
  OAI21X1 U2194 ( .A(n4497), .B(n2719), .C(n5625), .Y(n7829) );
  NAND2X1 U2195 ( .A(arr[1071]), .B(n2720), .Y(n5625) );
  OAI21X1 U2196 ( .A(n4499), .B(n2719), .C(n5626), .Y(n7830) );
  NAND2X1 U2197 ( .A(arr[1072]), .B(n2720), .Y(n5626) );
  OAI21X1 U2198 ( .A(n4501), .B(n2718), .C(n5627), .Y(n7831) );
  NAND2X1 U2199 ( .A(arr[1073]), .B(n2720), .Y(n5627) );
  OAI21X1 U2200 ( .A(n4503), .B(n2718), .C(n5628), .Y(n7832) );
  NAND2X1 U2201 ( .A(arr[1074]), .B(n2720), .Y(n5628) );
  OAI21X1 U2202 ( .A(n4505), .B(n2718), .C(n5629), .Y(n7833) );
  NAND2X1 U2203 ( .A(arr[1075]), .B(n2720), .Y(n5629) );
  OAI21X1 U2204 ( .A(n4507), .B(n2718), .C(n5630), .Y(n7834) );
  NAND2X1 U2205 ( .A(arr[1076]), .B(n2720), .Y(n5630) );
  OAI21X1 U2206 ( .A(n4509), .B(n2718), .C(n5631), .Y(n7835) );
  NAND2X1 U2207 ( .A(arr[1077]), .B(n2720), .Y(n5631) );
  OAI21X1 U2208 ( .A(n4511), .B(n2718), .C(n5632), .Y(n7836) );
  NAND2X1 U2209 ( .A(arr[1078]), .B(n2720), .Y(n5632) );
  OAI21X1 U2210 ( .A(n4513), .B(n2720), .C(n5633), .Y(n7837) );
  NAND2X1 U2211 ( .A(arr[1079]), .B(n2720), .Y(n5633) );
  OAI21X1 U2212 ( .A(n4515), .B(n2718), .C(n5634), .Y(n7838) );
  NAND2X1 U2213 ( .A(arr[1080]), .B(n2720), .Y(n5634) );
  OAI21X1 U2214 ( .A(n4517), .B(n2719), .C(n5635), .Y(n7839) );
  NAND2X1 U2215 ( .A(arr[1081]), .B(n2720), .Y(n5635) );
  OAI21X1 U2216 ( .A(n4519), .B(n2718), .C(n5636), .Y(n7840) );
  NAND2X1 U2217 ( .A(arr[1082]), .B(n2719), .Y(n5636) );
  OAI21X1 U2218 ( .A(n4521), .B(n2719), .C(n5637), .Y(n7841) );
  NAND2X1 U2219 ( .A(arr[1083]), .B(n2720), .Y(n5637) );
  OAI21X1 U2220 ( .A(n4523), .B(n2718), .C(n5638), .Y(n7842) );
  NAND2X1 U2221 ( .A(arr[1084]), .B(n2719), .Y(n5638) );
  OAI21X1 U2222 ( .A(n4525), .B(n2718), .C(n5639), .Y(n7843) );
  NAND2X1 U2223 ( .A(arr[1085]), .B(n2720), .Y(n5639) );
  OAI21X1 U2224 ( .A(n4527), .B(n2718), .C(n5640), .Y(n7844) );
  NAND2X1 U2225 ( .A(arr[1086]), .B(n2719), .Y(n5640) );
  OAI21X1 U2226 ( .A(n4529), .B(n2718), .C(n5641), .Y(n7845) );
  NAND2X1 U2227 ( .A(arr[1087]), .B(n2719), .Y(n5641) );
  OAI21X1 U2228 ( .A(n4531), .B(n2718), .C(n5642), .Y(n7846) );
  NAND2X1 U2229 ( .A(arr[1088]), .B(n2720), .Y(n5642) );
  OAI21X1 U2231 ( .A(n4467), .B(n2717), .C(n5645), .Y(n7847) );
  NAND2X1 U2232 ( .A(arr[1089]), .B(n2716), .Y(n5645) );
  OAI21X1 U2233 ( .A(n4469), .B(n2715), .C(n5646), .Y(n7848) );
  NAND2X1 U2234 ( .A(arr[1090]), .B(n2716), .Y(n5646) );
  OAI21X1 U2235 ( .A(n4471), .B(n2715), .C(n5647), .Y(n7849) );
  NAND2X1 U2236 ( .A(arr[1091]), .B(n2716), .Y(n5647) );
  OAI21X1 U2237 ( .A(n4473), .B(n2715), .C(n5648), .Y(n7850) );
  NAND2X1 U2238 ( .A(arr[1092]), .B(n2716), .Y(n5648) );
  OAI21X1 U2239 ( .A(n4475), .B(n2715), .C(n5649), .Y(n7851) );
  NAND2X1 U2240 ( .A(arr[1093]), .B(n2716), .Y(n5649) );
  OAI21X1 U2241 ( .A(n4477), .B(n2715), .C(n5650), .Y(n7852) );
  NAND2X1 U2242 ( .A(arr[1094]), .B(n2717), .Y(n5650) );
  OAI21X1 U2243 ( .A(n4479), .B(n2715), .C(n5651), .Y(n7853) );
  NAND2X1 U2244 ( .A(arr[1095]), .B(n2717), .Y(n5651) );
  OAI21X1 U2245 ( .A(n4481), .B(n2716), .C(n5652), .Y(n7854) );
  NAND2X1 U2246 ( .A(arr[1096]), .B(n2716), .Y(n5652) );
  OAI21X1 U2247 ( .A(n4483), .B(n2715), .C(n5653), .Y(n7855) );
  NAND2X1 U2248 ( .A(arr[1097]), .B(n2716), .Y(n5653) );
  OAI21X1 U2249 ( .A(n4485), .B(n2716), .C(n5654), .Y(n7856) );
  NAND2X1 U2250 ( .A(arr[1098]), .B(n2717), .Y(n5654) );
  OAI21X1 U2251 ( .A(n4487), .B(n2716), .C(n5655), .Y(n7857) );
  NAND2X1 U2252 ( .A(arr[1099]), .B(n2717), .Y(n5655) );
  OAI21X1 U2253 ( .A(n4489), .B(n2715), .C(n5656), .Y(n7858) );
  NAND2X1 U2254 ( .A(arr[1100]), .B(n2717), .Y(n5656) );
  OAI21X1 U2255 ( .A(n4491), .B(n2716), .C(n5657), .Y(n7859) );
  NAND2X1 U2256 ( .A(arr[1101]), .B(n2717), .Y(n5657) );
  OAI21X1 U2257 ( .A(n4493), .B(n2716), .C(n5658), .Y(n7860) );
  NAND2X1 U2258 ( .A(arr[1102]), .B(n2717), .Y(n5658) );
  OAI21X1 U2259 ( .A(n4495), .B(n2715), .C(n5659), .Y(n7861) );
  NAND2X1 U2260 ( .A(arr[1103]), .B(n2717), .Y(n5659) );
  OAI21X1 U2261 ( .A(n4497), .B(n2716), .C(n5660), .Y(n7862) );
  NAND2X1 U2262 ( .A(arr[1104]), .B(n2717), .Y(n5660) );
  OAI21X1 U2263 ( .A(n4499), .B(n2716), .C(n5661), .Y(n7863) );
  NAND2X1 U2264 ( .A(arr[1105]), .B(n2717), .Y(n5661) );
  OAI21X1 U2265 ( .A(n4501), .B(n2715), .C(n5662), .Y(n7864) );
  NAND2X1 U2266 ( .A(arr[1106]), .B(n2717), .Y(n5662) );
  OAI21X1 U2267 ( .A(n4503), .B(n2715), .C(n5663), .Y(n7865) );
  NAND2X1 U2268 ( .A(arr[1107]), .B(n2717), .Y(n5663) );
  OAI21X1 U2269 ( .A(n4505), .B(n2715), .C(n5664), .Y(n7866) );
  NAND2X1 U2270 ( .A(arr[1108]), .B(n2717), .Y(n5664) );
  OAI21X1 U2271 ( .A(n4507), .B(n2715), .C(n5665), .Y(n7867) );
  NAND2X1 U2272 ( .A(arr[1109]), .B(n2717), .Y(n5665) );
  OAI21X1 U2273 ( .A(n4509), .B(n2715), .C(n5666), .Y(n7868) );
  NAND2X1 U2274 ( .A(arr[1110]), .B(n2717), .Y(n5666) );
  OAI21X1 U2275 ( .A(n4511), .B(n2715), .C(n5667), .Y(n7869) );
  NAND2X1 U2276 ( .A(arr[1111]), .B(n2717), .Y(n5667) );
  OAI21X1 U2277 ( .A(n4513), .B(n2717), .C(n5668), .Y(n7870) );
  NAND2X1 U2278 ( .A(arr[1112]), .B(n2717), .Y(n5668) );
  OAI21X1 U2279 ( .A(n4515), .B(n2715), .C(n5669), .Y(n7871) );
  NAND2X1 U2280 ( .A(arr[1113]), .B(n2717), .Y(n5669) );
  OAI21X1 U2281 ( .A(n4517), .B(n2716), .C(n5670), .Y(n7872) );
  NAND2X1 U2282 ( .A(arr[1114]), .B(n2717), .Y(n5670) );
  OAI21X1 U2283 ( .A(n4519), .B(n2715), .C(n5671), .Y(n7873) );
  NAND2X1 U2284 ( .A(arr[1115]), .B(n2716), .Y(n5671) );
  OAI21X1 U2285 ( .A(n4521), .B(n2716), .C(n5672), .Y(n7874) );
  NAND2X1 U2286 ( .A(arr[1116]), .B(n2717), .Y(n5672) );
  OAI21X1 U2287 ( .A(n4523), .B(n2715), .C(n5673), .Y(n7875) );
  NAND2X1 U2288 ( .A(arr[1117]), .B(n2716), .Y(n5673) );
  OAI21X1 U2289 ( .A(n4525), .B(n2715), .C(n5674), .Y(n7876) );
  NAND2X1 U2290 ( .A(arr[1118]), .B(n2717), .Y(n5674) );
  OAI21X1 U2291 ( .A(n4527), .B(n2715), .C(n5675), .Y(n7877) );
  NAND2X1 U2292 ( .A(arr[1119]), .B(n2716), .Y(n5675) );
  OAI21X1 U2293 ( .A(n4529), .B(n2715), .C(n5676), .Y(n7878) );
  NAND2X1 U2294 ( .A(arr[1120]), .B(n2716), .Y(n5676) );
  OAI21X1 U2295 ( .A(n4531), .B(n2715), .C(n5677), .Y(n7879) );
  NAND2X1 U2296 ( .A(arr[1121]), .B(n2717), .Y(n5677) );
  AND2X1 U2298 ( .A(n5679), .B(n5680), .Y(n4534) );
  OAI21X1 U2299 ( .A(n4467), .B(n2714), .C(n5682), .Y(n7880) );
  NAND2X1 U2300 ( .A(arr[1122]), .B(n2713), .Y(n5682) );
  OAI21X1 U2301 ( .A(n4469), .B(n2712), .C(n5683), .Y(n7881) );
  NAND2X1 U2302 ( .A(arr[1123]), .B(n2713), .Y(n5683) );
  OAI21X1 U2303 ( .A(n4471), .B(n2712), .C(n5684), .Y(n7882) );
  NAND2X1 U2304 ( .A(arr[1124]), .B(n2713), .Y(n5684) );
  OAI21X1 U2305 ( .A(n4473), .B(n2712), .C(n5685), .Y(n7883) );
  NAND2X1 U2306 ( .A(arr[1125]), .B(n2713), .Y(n5685) );
  OAI21X1 U2307 ( .A(n4475), .B(n2712), .C(n5686), .Y(n7884) );
  NAND2X1 U2308 ( .A(arr[1126]), .B(n2713), .Y(n5686) );
  OAI21X1 U2309 ( .A(n4477), .B(n2712), .C(n5687), .Y(n7885) );
  NAND2X1 U2310 ( .A(arr[1127]), .B(n2714), .Y(n5687) );
  OAI21X1 U2311 ( .A(n4479), .B(n2712), .C(n5688), .Y(n7886) );
  NAND2X1 U2312 ( .A(arr[1128]), .B(n2714), .Y(n5688) );
  OAI21X1 U2313 ( .A(n4481), .B(n2713), .C(n5689), .Y(n7887) );
  NAND2X1 U2314 ( .A(arr[1129]), .B(n2713), .Y(n5689) );
  OAI21X1 U2315 ( .A(n4483), .B(n2712), .C(n5690), .Y(n7888) );
  NAND2X1 U2316 ( .A(arr[1130]), .B(n2713), .Y(n5690) );
  OAI21X1 U2317 ( .A(n4485), .B(n2713), .C(n5691), .Y(n7889) );
  NAND2X1 U2318 ( .A(arr[1131]), .B(n2714), .Y(n5691) );
  OAI21X1 U2319 ( .A(n4487), .B(n2713), .C(n5692), .Y(n7890) );
  NAND2X1 U2320 ( .A(arr[1132]), .B(n2714), .Y(n5692) );
  OAI21X1 U2321 ( .A(n4489), .B(n2712), .C(n5693), .Y(n7891) );
  NAND2X1 U2322 ( .A(arr[1133]), .B(n2714), .Y(n5693) );
  OAI21X1 U2323 ( .A(n4491), .B(n2713), .C(n5694), .Y(n7892) );
  NAND2X1 U2324 ( .A(arr[1134]), .B(n2714), .Y(n5694) );
  OAI21X1 U2325 ( .A(n4493), .B(n2713), .C(n5695), .Y(n7893) );
  NAND2X1 U2326 ( .A(arr[1135]), .B(n2714), .Y(n5695) );
  OAI21X1 U2327 ( .A(n4495), .B(n2712), .C(n5696), .Y(n7894) );
  NAND2X1 U2328 ( .A(arr[1136]), .B(n2714), .Y(n5696) );
  OAI21X1 U2329 ( .A(n4497), .B(n2713), .C(n5697), .Y(n7895) );
  NAND2X1 U2330 ( .A(arr[1137]), .B(n2714), .Y(n5697) );
  OAI21X1 U2331 ( .A(n4499), .B(n2713), .C(n5698), .Y(n7896) );
  NAND2X1 U2332 ( .A(arr[1138]), .B(n2714), .Y(n5698) );
  OAI21X1 U2333 ( .A(n4501), .B(n2712), .C(n5699), .Y(n7897) );
  NAND2X1 U2334 ( .A(arr[1139]), .B(n2714), .Y(n5699) );
  OAI21X1 U2335 ( .A(n4503), .B(n2712), .C(n5700), .Y(n7898) );
  NAND2X1 U2336 ( .A(arr[1140]), .B(n2714), .Y(n5700) );
  OAI21X1 U2337 ( .A(n4505), .B(n2712), .C(n5701), .Y(n7899) );
  NAND2X1 U2338 ( .A(arr[1141]), .B(n2714), .Y(n5701) );
  OAI21X1 U2339 ( .A(n4507), .B(n2712), .C(n5702), .Y(n7900) );
  NAND2X1 U2340 ( .A(arr[1142]), .B(n2714), .Y(n5702) );
  OAI21X1 U2341 ( .A(n4509), .B(n2712), .C(n5703), .Y(n7901) );
  NAND2X1 U2342 ( .A(arr[1143]), .B(n2714), .Y(n5703) );
  OAI21X1 U2343 ( .A(n4511), .B(n2712), .C(n5704), .Y(n7902) );
  NAND2X1 U2344 ( .A(arr[1144]), .B(n2714), .Y(n5704) );
  OAI21X1 U2345 ( .A(n4513), .B(n2714), .C(n5705), .Y(n7903) );
  NAND2X1 U2346 ( .A(arr[1145]), .B(n2714), .Y(n5705) );
  OAI21X1 U2347 ( .A(n4515), .B(n2712), .C(n5706), .Y(n7904) );
  NAND2X1 U2348 ( .A(arr[1146]), .B(n2714), .Y(n5706) );
  OAI21X1 U2349 ( .A(n4517), .B(n2713), .C(n5707), .Y(n7905) );
  NAND2X1 U2350 ( .A(arr[1147]), .B(n2714), .Y(n5707) );
  OAI21X1 U2351 ( .A(n4519), .B(n2712), .C(n5708), .Y(n7906) );
  NAND2X1 U2352 ( .A(arr[1148]), .B(n2713), .Y(n5708) );
  OAI21X1 U2353 ( .A(n4521), .B(n2713), .C(n5709), .Y(n7907) );
  NAND2X1 U2354 ( .A(arr[1149]), .B(n2714), .Y(n5709) );
  OAI21X1 U2355 ( .A(n4523), .B(n2712), .C(n5710), .Y(n7908) );
  NAND2X1 U2356 ( .A(arr[1150]), .B(n2713), .Y(n5710) );
  OAI21X1 U2357 ( .A(n4525), .B(n2712), .C(n5711), .Y(n7909) );
  NAND2X1 U2358 ( .A(arr[1151]), .B(n2714), .Y(n5711) );
  OAI21X1 U2359 ( .A(n4527), .B(n2712), .C(n5712), .Y(n7910) );
  NAND2X1 U2360 ( .A(arr[1152]), .B(n2713), .Y(n5712) );
  OAI21X1 U2361 ( .A(n4529), .B(n2712), .C(n5713), .Y(n7911) );
  NAND2X1 U2362 ( .A(arr[1153]), .B(n2713), .Y(n5713) );
  OAI21X1 U2363 ( .A(n4531), .B(n2712), .C(n5714), .Y(n7912) );
  NAND2X1 U2364 ( .A(arr[1154]), .B(n2714), .Y(n5714) );
  OAI21X1 U2366 ( .A(n4467), .B(n2711), .C(n5716), .Y(n7913) );
  NAND2X1 U2367 ( .A(arr[1155]), .B(n2710), .Y(n5716) );
  OAI21X1 U2368 ( .A(n4469), .B(n2709), .C(n5717), .Y(n7914) );
  NAND2X1 U2369 ( .A(arr[1156]), .B(n2710), .Y(n5717) );
  OAI21X1 U2370 ( .A(n4471), .B(n2709), .C(n5718), .Y(n7915) );
  NAND2X1 U2371 ( .A(arr[1157]), .B(n2710), .Y(n5718) );
  OAI21X1 U2372 ( .A(n4473), .B(n2709), .C(n5719), .Y(n7916) );
  NAND2X1 U2373 ( .A(arr[1158]), .B(n2710), .Y(n5719) );
  OAI21X1 U2374 ( .A(n4475), .B(n2709), .C(n5720), .Y(n7917) );
  NAND2X1 U2375 ( .A(arr[1159]), .B(n2710), .Y(n5720) );
  OAI21X1 U2376 ( .A(n4477), .B(n2709), .C(n5721), .Y(n7918) );
  NAND2X1 U2377 ( .A(arr[1160]), .B(n2711), .Y(n5721) );
  OAI21X1 U2378 ( .A(n4479), .B(n2709), .C(n5722), .Y(n7919) );
  NAND2X1 U2379 ( .A(arr[1161]), .B(n2711), .Y(n5722) );
  OAI21X1 U2380 ( .A(n4481), .B(n2710), .C(n5723), .Y(n7920) );
  NAND2X1 U2381 ( .A(arr[1162]), .B(n2710), .Y(n5723) );
  OAI21X1 U2382 ( .A(n4483), .B(n2709), .C(n5724), .Y(n7921) );
  NAND2X1 U2383 ( .A(arr[1163]), .B(n2710), .Y(n5724) );
  OAI21X1 U2384 ( .A(n4485), .B(n2710), .C(n5725), .Y(n7922) );
  NAND2X1 U2385 ( .A(arr[1164]), .B(n2711), .Y(n5725) );
  OAI21X1 U2386 ( .A(n4487), .B(n2710), .C(n5726), .Y(n7923) );
  NAND2X1 U2387 ( .A(arr[1165]), .B(n2711), .Y(n5726) );
  OAI21X1 U2388 ( .A(n4489), .B(n2709), .C(n5727), .Y(n7924) );
  NAND2X1 U2389 ( .A(arr[1166]), .B(n2711), .Y(n5727) );
  OAI21X1 U2390 ( .A(n4491), .B(n2710), .C(n5728), .Y(n7925) );
  NAND2X1 U2391 ( .A(arr[1167]), .B(n2711), .Y(n5728) );
  OAI21X1 U2392 ( .A(n4493), .B(n2710), .C(n5729), .Y(n7926) );
  NAND2X1 U2393 ( .A(arr[1168]), .B(n2711), .Y(n5729) );
  OAI21X1 U2394 ( .A(n4495), .B(n2709), .C(n5730), .Y(n7927) );
  NAND2X1 U2395 ( .A(arr[1169]), .B(n2711), .Y(n5730) );
  OAI21X1 U2396 ( .A(n4497), .B(n2710), .C(n5731), .Y(n7928) );
  NAND2X1 U2397 ( .A(arr[1170]), .B(n2711), .Y(n5731) );
  OAI21X1 U2398 ( .A(n4499), .B(n2710), .C(n5732), .Y(n7929) );
  NAND2X1 U2399 ( .A(arr[1171]), .B(n2711), .Y(n5732) );
  OAI21X1 U2400 ( .A(n4501), .B(n2709), .C(n5733), .Y(n7930) );
  NAND2X1 U2401 ( .A(arr[1172]), .B(n2711), .Y(n5733) );
  OAI21X1 U2402 ( .A(n4503), .B(n2709), .C(n5734), .Y(n7931) );
  NAND2X1 U2403 ( .A(arr[1173]), .B(n2711), .Y(n5734) );
  OAI21X1 U2404 ( .A(n4505), .B(n2709), .C(n5735), .Y(n7932) );
  NAND2X1 U2405 ( .A(arr[1174]), .B(n2711), .Y(n5735) );
  OAI21X1 U2406 ( .A(n4507), .B(n2709), .C(n5736), .Y(n7933) );
  NAND2X1 U2407 ( .A(arr[1175]), .B(n2711), .Y(n5736) );
  OAI21X1 U2408 ( .A(n4509), .B(n2709), .C(n5737), .Y(n7934) );
  NAND2X1 U2409 ( .A(arr[1176]), .B(n2711), .Y(n5737) );
  OAI21X1 U2410 ( .A(n4511), .B(n2709), .C(n5738), .Y(n7935) );
  NAND2X1 U2411 ( .A(arr[1177]), .B(n2711), .Y(n5738) );
  OAI21X1 U2412 ( .A(n4513), .B(n2711), .C(n5739), .Y(n7936) );
  NAND2X1 U2413 ( .A(arr[1178]), .B(n2711), .Y(n5739) );
  OAI21X1 U2414 ( .A(n4515), .B(n2709), .C(n5740), .Y(n7937) );
  NAND2X1 U2415 ( .A(arr[1179]), .B(n2711), .Y(n5740) );
  OAI21X1 U2416 ( .A(n4517), .B(n2710), .C(n5741), .Y(n7938) );
  NAND2X1 U2417 ( .A(arr[1180]), .B(n2711), .Y(n5741) );
  OAI21X1 U2418 ( .A(n4519), .B(n2709), .C(n5742), .Y(n7939) );
  NAND2X1 U2419 ( .A(arr[1181]), .B(n2710), .Y(n5742) );
  OAI21X1 U2420 ( .A(n4521), .B(n2710), .C(n5743), .Y(n7940) );
  NAND2X1 U2421 ( .A(arr[1182]), .B(n2711), .Y(n5743) );
  OAI21X1 U2422 ( .A(n4523), .B(n2709), .C(n5744), .Y(n7941) );
  NAND2X1 U2423 ( .A(arr[1183]), .B(n2710), .Y(n5744) );
  OAI21X1 U2424 ( .A(n4525), .B(n2709), .C(n5745), .Y(n7942) );
  NAND2X1 U2425 ( .A(arr[1184]), .B(n2711), .Y(n5745) );
  OAI21X1 U2426 ( .A(n4527), .B(n2709), .C(n5746), .Y(n7943) );
  NAND2X1 U2427 ( .A(arr[1185]), .B(n2710), .Y(n5746) );
  OAI21X1 U2428 ( .A(n4529), .B(n2709), .C(n5747), .Y(n7944) );
  NAND2X1 U2429 ( .A(arr[1186]), .B(n2710), .Y(n5747) );
  OAI21X1 U2430 ( .A(n4531), .B(n2709), .C(n5748), .Y(n7945) );
  NAND2X1 U2431 ( .A(arr[1187]), .B(n2711), .Y(n5748) );
  AND2X1 U2433 ( .A(n5749), .B(n5679), .Y(n4604) );
  OAI21X1 U2434 ( .A(n4467), .B(n2708), .C(n5751), .Y(n7946) );
  NAND2X1 U2435 ( .A(arr[1188]), .B(n2707), .Y(n5751) );
  OAI21X1 U2436 ( .A(n4469), .B(n2706), .C(n5752), .Y(n7947) );
  NAND2X1 U2437 ( .A(arr[1189]), .B(n2707), .Y(n5752) );
  OAI21X1 U2438 ( .A(n4471), .B(n2706), .C(n5753), .Y(n7948) );
  NAND2X1 U2439 ( .A(arr[1190]), .B(n2707), .Y(n5753) );
  OAI21X1 U2440 ( .A(n4473), .B(n2706), .C(n5754), .Y(n7949) );
  NAND2X1 U2441 ( .A(arr[1191]), .B(n2707), .Y(n5754) );
  OAI21X1 U2442 ( .A(n4475), .B(n2706), .C(n5755), .Y(n7950) );
  NAND2X1 U2443 ( .A(arr[1192]), .B(n2707), .Y(n5755) );
  OAI21X1 U2444 ( .A(n4477), .B(n2706), .C(n5756), .Y(n7951) );
  NAND2X1 U2445 ( .A(arr[1193]), .B(n2708), .Y(n5756) );
  OAI21X1 U2446 ( .A(n4479), .B(n2706), .C(n5757), .Y(n7952) );
  NAND2X1 U2447 ( .A(arr[1194]), .B(n2708), .Y(n5757) );
  OAI21X1 U2448 ( .A(n4481), .B(n2707), .C(n5758), .Y(n7953) );
  NAND2X1 U2449 ( .A(arr[1195]), .B(n2707), .Y(n5758) );
  OAI21X1 U2450 ( .A(n4483), .B(n2706), .C(n5759), .Y(n7954) );
  NAND2X1 U2451 ( .A(arr[1196]), .B(n2707), .Y(n5759) );
  OAI21X1 U2452 ( .A(n4485), .B(n2707), .C(n5760), .Y(n7955) );
  NAND2X1 U2453 ( .A(arr[1197]), .B(n2708), .Y(n5760) );
  OAI21X1 U2454 ( .A(n4487), .B(n2707), .C(n5761), .Y(n7956) );
  NAND2X1 U2455 ( .A(arr[1198]), .B(n2708), .Y(n5761) );
  OAI21X1 U2456 ( .A(n4489), .B(n2706), .C(n5762), .Y(n7957) );
  NAND2X1 U2457 ( .A(arr[1199]), .B(n2708), .Y(n5762) );
  OAI21X1 U2458 ( .A(n4491), .B(n2707), .C(n5763), .Y(n7958) );
  NAND2X1 U2459 ( .A(arr[1200]), .B(n2708), .Y(n5763) );
  OAI21X1 U2460 ( .A(n4493), .B(n2707), .C(n5764), .Y(n7959) );
  NAND2X1 U2461 ( .A(arr[1201]), .B(n2708), .Y(n5764) );
  OAI21X1 U2462 ( .A(n4495), .B(n2706), .C(n5765), .Y(n7960) );
  NAND2X1 U2463 ( .A(arr[1202]), .B(n2708), .Y(n5765) );
  OAI21X1 U2464 ( .A(n4497), .B(n2707), .C(n5766), .Y(n7961) );
  NAND2X1 U2465 ( .A(arr[1203]), .B(n2708), .Y(n5766) );
  OAI21X1 U2466 ( .A(n4499), .B(n2707), .C(n5767), .Y(n7962) );
  NAND2X1 U2467 ( .A(arr[1204]), .B(n2708), .Y(n5767) );
  OAI21X1 U2468 ( .A(n4501), .B(n2706), .C(n5768), .Y(n7963) );
  NAND2X1 U2469 ( .A(arr[1205]), .B(n2708), .Y(n5768) );
  OAI21X1 U2470 ( .A(n4503), .B(n2706), .C(n5769), .Y(n7964) );
  NAND2X1 U2471 ( .A(arr[1206]), .B(n2708), .Y(n5769) );
  OAI21X1 U2472 ( .A(n4505), .B(n2706), .C(n5770), .Y(n7965) );
  NAND2X1 U2473 ( .A(arr[1207]), .B(n2708), .Y(n5770) );
  OAI21X1 U2474 ( .A(n4507), .B(n2706), .C(n5771), .Y(n7966) );
  NAND2X1 U2475 ( .A(arr[1208]), .B(n2708), .Y(n5771) );
  OAI21X1 U2476 ( .A(n4509), .B(n2706), .C(n5772), .Y(n7967) );
  NAND2X1 U2477 ( .A(arr[1209]), .B(n2708), .Y(n5772) );
  OAI21X1 U2478 ( .A(n4511), .B(n2706), .C(n5773), .Y(n7968) );
  NAND2X1 U2479 ( .A(arr[1210]), .B(n2708), .Y(n5773) );
  OAI21X1 U2480 ( .A(n4513), .B(n2708), .C(n5774), .Y(n7969) );
  NAND2X1 U2481 ( .A(arr[1211]), .B(n2708), .Y(n5774) );
  OAI21X1 U2482 ( .A(n4515), .B(n2706), .C(n5775), .Y(n7970) );
  NAND2X1 U2483 ( .A(arr[1212]), .B(n2708), .Y(n5775) );
  OAI21X1 U2484 ( .A(n4517), .B(n2707), .C(n5776), .Y(n7971) );
  NAND2X1 U2485 ( .A(arr[1213]), .B(n2708), .Y(n5776) );
  OAI21X1 U2486 ( .A(n4519), .B(n2706), .C(n5777), .Y(n7972) );
  NAND2X1 U2487 ( .A(arr[1214]), .B(n2707), .Y(n5777) );
  OAI21X1 U2488 ( .A(n4521), .B(n2707), .C(n5778), .Y(n7973) );
  NAND2X1 U2489 ( .A(arr[1215]), .B(n2708), .Y(n5778) );
  OAI21X1 U2490 ( .A(n4523), .B(n2706), .C(n5779), .Y(n7974) );
  NAND2X1 U2491 ( .A(arr[1216]), .B(n2707), .Y(n5779) );
  OAI21X1 U2492 ( .A(n4525), .B(n2706), .C(n5780), .Y(n7975) );
  NAND2X1 U2493 ( .A(arr[1217]), .B(n2708), .Y(n5780) );
  OAI21X1 U2494 ( .A(n4527), .B(n2706), .C(n5781), .Y(n7976) );
  NAND2X1 U2495 ( .A(arr[1218]), .B(n2707), .Y(n5781) );
  OAI21X1 U2496 ( .A(n4529), .B(n2706), .C(n5782), .Y(n7977) );
  NAND2X1 U2497 ( .A(arr[1219]), .B(n2707), .Y(n5782) );
  OAI21X1 U2498 ( .A(n4531), .B(n2706), .C(n5783), .Y(n7978) );
  NAND2X1 U2499 ( .A(arr[1220]), .B(n2708), .Y(n5783) );
  OAI21X1 U2501 ( .A(n4467), .B(n2705), .C(n5785), .Y(n7979) );
  NAND2X1 U2502 ( .A(arr[1221]), .B(n2704), .Y(n5785) );
  OAI21X1 U2503 ( .A(n4469), .B(n2703), .C(n5786), .Y(n7980) );
  NAND2X1 U2504 ( .A(arr[1222]), .B(n2704), .Y(n5786) );
  OAI21X1 U2505 ( .A(n4471), .B(n2703), .C(n5787), .Y(n7981) );
  NAND2X1 U2506 ( .A(arr[1223]), .B(n2704), .Y(n5787) );
  OAI21X1 U2507 ( .A(n4473), .B(n2703), .C(n5788), .Y(n7982) );
  NAND2X1 U2508 ( .A(arr[1224]), .B(n2704), .Y(n5788) );
  OAI21X1 U2509 ( .A(n4475), .B(n2703), .C(n5789), .Y(n7983) );
  NAND2X1 U2510 ( .A(arr[1225]), .B(n2704), .Y(n5789) );
  OAI21X1 U2511 ( .A(n4477), .B(n2703), .C(n5790), .Y(n7984) );
  NAND2X1 U2512 ( .A(arr[1226]), .B(n2705), .Y(n5790) );
  OAI21X1 U2513 ( .A(n4479), .B(n2703), .C(n5791), .Y(n7985) );
  NAND2X1 U2514 ( .A(arr[1227]), .B(n2705), .Y(n5791) );
  OAI21X1 U2515 ( .A(n4481), .B(n2704), .C(n5792), .Y(n7986) );
  NAND2X1 U2516 ( .A(arr[1228]), .B(n2704), .Y(n5792) );
  OAI21X1 U2517 ( .A(n4483), .B(n2703), .C(n5793), .Y(n7987) );
  NAND2X1 U2518 ( .A(arr[1229]), .B(n2704), .Y(n5793) );
  OAI21X1 U2519 ( .A(n4485), .B(n2704), .C(n5794), .Y(n7988) );
  NAND2X1 U2520 ( .A(arr[1230]), .B(n2705), .Y(n5794) );
  OAI21X1 U2521 ( .A(n4487), .B(n2704), .C(n5795), .Y(n7989) );
  NAND2X1 U2522 ( .A(arr[1231]), .B(n2705), .Y(n5795) );
  OAI21X1 U2523 ( .A(n4489), .B(n2703), .C(n5796), .Y(n7990) );
  NAND2X1 U2524 ( .A(arr[1232]), .B(n2705), .Y(n5796) );
  OAI21X1 U2525 ( .A(n4491), .B(n2704), .C(n5797), .Y(n7991) );
  NAND2X1 U2526 ( .A(arr[1233]), .B(n2705), .Y(n5797) );
  OAI21X1 U2527 ( .A(n4493), .B(n2704), .C(n5798), .Y(n7992) );
  NAND2X1 U2528 ( .A(arr[1234]), .B(n2705), .Y(n5798) );
  OAI21X1 U2529 ( .A(n4495), .B(n2703), .C(n5799), .Y(n7993) );
  NAND2X1 U2530 ( .A(arr[1235]), .B(n2705), .Y(n5799) );
  OAI21X1 U2531 ( .A(n4497), .B(n2704), .C(n5800), .Y(n7994) );
  NAND2X1 U2532 ( .A(arr[1236]), .B(n2705), .Y(n5800) );
  OAI21X1 U2533 ( .A(n4499), .B(n2704), .C(n5801), .Y(n7995) );
  NAND2X1 U2534 ( .A(arr[1237]), .B(n2705), .Y(n5801) );
  OAI21X1 U2535 ( .A(n4501), .B(n2703), .C(n5802), .Y(n7996) );
  NAND2X1 U2536 ( .A(arr[1238]), .B(n2705), .Y(n5802) );
  OAI21X1 U2537 ( .A(n4503), .B(n2703), .C(n5803), .Y(n7997) );
  NAND2X1 U2538 ( .A(arr[1239]), .B(n2705), .Y(n5803) );
  OAI21X1 U2539 ( .A(n4505), .B(n2703), .C(n5804), .Y(n7998) );
  NAND2X1 U2540 ( .A(arr[1240]), .B(n2705), .Y(n5804) );
  OAI21X1 U2541 ( .A(n4507), .B(n2703), .C(n5805), .Y(n7999) );
  NAND2X1 U2542 ( .A(arr[1241]), .B(n2705), .Y(n5805) );
  OAI21X1 U2543 ( .A(n4509), .B(n2703), .C(n5806), .Y(n8000) );
  NAND2X1 U2544 ( .A(arr[1242]), .B(n2705), .Y(n5806) );
  OAI21X1 U2545 ( .A(n4511), .B(n2703), .C(n5807), .Y(n8001) );
  NAND2X1 U2546 ( .A(arr[1243]), .B(n2705), .Y(n5807) );
  OAI21X1 U2547 ( .A(n4513), .B(n2705), .C(n5808), .Y(n8002) );
  NAND2X1 U2548 ( .A(arr[1244]), .B(n2705), .Y(n5808) );
  OAI21X1 U2549 ( .A(n4515), .B(n2703), .C(n5809), .Y(n8003) );
  NAND2X1 U2550 ( .A(arr[1245]), .B(n2705), .Y(n5809) );
  OAI21X1 U2551 ( .A(n4517), .B(n2704), .C(n5810), .Y(n8004) );
  NAND2X1 U2552 ( .A(arr[1246]), .B(n2705), .Y(n5810) );
  OAI21X1 U2553 ( .A(n4519), .B(n2703), .C(n5811), .Y(n8005) );
  NAND2X1 U2554 ( .A(arr[1247]), .B(n2704), .Y(n5811) );
  OAI21X1 U2555 ( .A(n4521), .B(n2704), .C(n5812), .Y(n8006) );
  NAND2X1 U2556 ( .A(arr[1248]), .B(n2705), .Y(n5812) );
  OAI21X1 U2557 ( .A(n4523), .B(n2703), .C(n5813), .Y(n8007) );
  NAND2X1 U2558 ( .A(arr[1249]), .B(n2704), .Y(n5813) );
  OAI21X1 U2559 ( .A(n4525), .B(n2703), .C(n5814), .Y(n8008) );
  NAND2X1 U2560 ( .A(arr[1250]), .B(n2705), .Y(n5814) );
  OAI21X1 U2561 ( .A(n4527), .B(n2703), .C(n5815), .Y(n8009) );
  NAND2X1 U2562 ( .A(arr[1251]), .B(n2704), .Y(n5815) );
  OAI21X1 U2563 ( .A(n4529), .B(n2703), .C(n5816), .Y(n8010) );
  NAND2X1 U2564 ( .A(arr[1252]), .B(n2704), .Y(n5816) );
  OAI21X1 U2565 ( .A(n4531), .B(n2703), .C(n5817), .Y(n8011) );
  NAND2X1 U2566 ( .A(arr[1253]), .B(n2705), .Y(n5817) );
  AND2X1 U2568 ( .A(n5818), .B(n5679), .Y(n4673) );
  OAI21X1 U2569 ( .A(n4467), .B(n2702), .C(n5820), .Y(n8012) );
  NAND2X1 U2570 ( .A(arr[1254]), .B(n2701), .Y(n5820) );
  OAI21X1 U2571 ( .A(n4469), .B(n2700), .C(n5821), .Y(n8013) );
  NAND2X1 U2572 ( .A(arr[1255]), .B(n2701), .Y(n5821) );
  OAI21X1 U2573 ( .A(n4471), .B(n2700), .C(n5822), .Y(n8014) );
  NAND2X1 U2574 ( .A(arr[1256]), .B(n2701), .Y(n5822) );
  OAI21X1 U2575 ( .A(n4473), .B(n2700), .C(n5823), .Y(n8015) );
  NAND2X1 U2576 ( .A(arr[1257]), .B(n2701), .Y(n5823) );
  OAI21X1 U2577 ( .A(n4475), .B(n2700), .C(n5824), .Y(n8016) );
  NAND2X1 U2578 ( .A(arr[1258]), .B(n2701), .Y(n5824) );
  OAI21X1 U2579 ( .A(n4477), .B(n2700), .C(n5825), .Y(n8017) );
  NAND2X1 U2580 ( .A(arr[1259]), .B(n2702), .Y(n5825) );
  OAI21X1 U2581 ( .A(n4479), .B(n2700), .C(n5826), .Y(n8018) );
  NAND2X1 U2582 ( .A(arr[1260]), .B(n2702), .Y(n5826) );
  OAI21X1 U2583 ( .A(n4481), .B(n2701), .C(n5827), .Y(n8019) );
  NAND2X1 U2584 ( .A(arr[1261]), .B(n2701), .Y(n5827) );
  OAI21X1 U2585 ( .A(n4483), .B(n2700), .C(n5828), .Y(n8020) );
  NAND2X1 U2586 ( .A(arr[1262]), .B(n2701), .Y(n5828) );
  OAI21X1 U2587 ( .A(n4485), .B(n2701), .C(n5829), .Y(n8021) );
  NAND2X1 U2588 ( .A(arr[1263]), .B(n2702), .Y(n5829) );
  OAI21X1 U2589 ( .A(n4487), .B(n2701), .C(n5830), .Y(n8022) );
  NAND2X1 U2590 ( .A(arr[1264]), .B(n2702), .Y(n5830) );
  OAI21X1 U2591 ( .A(n4489), .B(n2700), .C(n5831), .Y(n8023) );
  NAND2X1 U2592 ( .A(arr[1265]), .B(n2702), .Y(n5831) );
  OAI21X1 U2593 ( .A(n4491), .B(n2701), .C(n5832), .Y(n8024) );
  NAND2X1 U2594 ( .A(arr[1266]), .B(n2702), .Y(n5832) );
  OAI21X1 U2595 ( .A(n4493), .B(n2701), .C(n5833), .Y(n8025) );
  NAND2X1 U2596 ( .A(arr[1267]), .B(n2702), .Y(n5833) );
  OAI21X1 U2597 ( .A(n4495), .B(n2700), .C(n5834), .Y(n8026) );
  NAND2X1 U2598 ( .A(arr[1268]), .B(n2702), .Y(n5834) );
  OAI21X1 U2599 ( .A(n4497), .B(n2701), .C(n5835), .Y(n8027) );
  NAND2X1 U2600 ( .A(arr[1269]), .B(n2702), .Y(n5835) );
  OAI21X1 U2601 ( .A(n4499), .B(n2701), .C(n5836), .Y(n8028) );
  NAND2X1 U2602 ( .A(arr[1270]), .B(n2702), .Y(n5836) );
  OAI21X1 U2603 ( .A(n4501), .B(n2700), .C(n5837), .Y(n8029) );
  NAND2X1 U2604 ( .A(arr[1271]), .B(n2702), .Y(n5837) );
  OAI21X1 U2605 ( .A(n4503), .B(n2700), .C(n5838), .Y(n8030) );
  NAND2X1 U2606 ( .A(arr[1272]), .B(n2702), .Y(n5838) );
  OAI21X1 U2607 ( .A(n4505), .B(n2700), .C(n5839), .Y(n8031) );
  NAND2X1 U2608 ( .A(arr[1273]), .B(n2702), .Y(n5839) );
  OAI21X1 U2609 ( .A(n4507), .B(n2700), .C(n5840), .Y(n8032) );
  NAND2X1 U2610 ( .A(arr[1274]), .B(n2702), .Y(n5840) );
  OAI21X1 U2611 ( .A(n4509), .B(n2700), .C(n5841), .Y(n8033) );
  NAND2X1 U2612 ( .A(arr[1275]), .B(n2702), .Y(n5841) );
  OAI21X1 U2613 ( .A(n4511), .B(n2700), .C(n5842), .Y(n8034) );
  NAND2X1 U2614 ( .A(arr[1276]), .B(n2702), .Y(n5842) );
  OAI21X1 U2615 ( .A(n4513), .B(n2702), .C(n5843), .Y(n8035) );
  NAND2X1 U2616 ( .A(arr[1277]), .B(n2702), .Y(n5843) );
  OAI21X1 U2617 ( .A(n4515), .B(n2700), .C(n5844), .Y(n8036) );
  NAND2X1 U2618 ( .A(arr[1278]), .B(n2702), .Y(n5844) );
  OAI21X1 U2619 ( .A(n4517), .B(n2701), .C(n5845), .Y(n8037) );
  NAND2X1 U2620 ( .A(arr[1279]), .B(n2702), .Y(n5845) );
  OAI21X1 U2621 ( .A(n4519), .B(n2700), .C(n5846), .Y(n8038) );
  NAND2X1 U2622 ( .A(arr[1280]), .B(n2701), .Y(n5846) );
  OAI21X1 U2623 ( .A(n4521), .B(n2701), .C(n5847), .Y(n8039) );
  NAND2X1 U2624 ( .A(arr[1281]), .B(n2702), .Y(n5847) );
  OAI21X1 U2625 ( .A(n4523), .B(n2700), .C(n5848), .Y(n8040) );
  NAND2X1 U2626 ( .A(arr[1282]), .B(n2701), .Y(n5848) );
  OAI21X1 U2627 ( .A(n4525), .B(n2700), .C(n5849), .Y(n8041) );
  NAND2X1 U2628 ( .A(arr[1283]), .B(n2702), .Y(n5849) );
  OAI21X1 U2629 ( .A(n4527), .B(n2700), .C(n5850), .Y(n8042) );
  NAND2X1 U2630 ( .A(arr[1284]), .B(n2701), .Y(n5850) );
  OAI21X1 U2631 ( .A(n4529), .B(n2700), .C(n5851), .Y(n8043) );
  NAND2X1 U2632 ( .A(arr[1285]), .B(n2701), .Y(n5851) );
  OAI21X1 U2633 ( .A(n4531), .B(n2700), .C(n5852), .Y(n8044) );
  NAND2X1 U2634 ( .A(arr[1286]), .B(n2702), .Y(n5852) );
  OAI21X1 U2636 ( .A(n4467), .B(n2699), .C(n5854), .Y(n8045) );
  NAND2X1 U2637 ( .A(arr[1287]), .B(n2698), .Y(n5854) );
  OAI21X1 U2638 ( .A(n4469), .B(n2697), .C(n5855), .Y(n8046) );
  NAND2X1 U2639 ( .A(arr[1288]), .B(n2698), .Y(n5855) );
  OAI21X1 U2640 ( .A(n4471), .B(n2697), .C(n5856), .Y(n8047) );
  NAND2X1 U2641 ( .A(arr[1289]), .B(n2698), .Y(n5856) );
  OAI21X1 U2642 ( .A(n4473), .B(n2697), .C(n5857), .Y(n8048) );
  NAND2X1 U2643 ( .A(arr[1290]), .B(n2698), .Y(n5857) );
  OAI21X1 U2644 ( .A(n4475), .B(n2697), .C(n5858), .Y(n8049) );
  NAND2X1 U2645 ( .A(arr[1291]), .B(n2698), .Y(n5858) );
  OAI21X1 U2646 ( .A(n4477), .B(n2697), .C(n5859), .Y(n8050) );
  NAND2X1 U2647 ( .A(arr[1292]), .B(n2699), .Y(n5859) );
  OAI21X1 U2648 ( .A(n4479), .B(n2697), .C(n5860), .Y(n8051) );
  NAND2X1 U2649 ( .A(arr[1293]), .B(n2699), .Y(n5860) );
  OAI21X1 U2650 ( .A(n4481), .B(n2698), .C(n5861), .Y(n8052) );
  NAND2X1 U2651 ( .A(arr[1294]), .B(n2698), .Y(n5861) );
  OAI21X1 U2652 ( .A(n4483), .B(n2697), .C(n5862), .Y(n8053) );
  NAND2X1 U2653 ( .A(arr[1295]), .B(n2698), .Y(n5862) );
  OAI21X1 U2654 ( .A(n4485), .B(n2698), .C(n5863), .Y(n8054) );
  NAND2X1 U2655 ( .A(arr[1296]), .B(n2699), .Y(n5863) );
  OAI21X1 U2656 ( .A(n4487), .B(n2698), .C(n5864), .Y(n8055) );
  NAND2X1 U2657 ( .A(arr[1297]), .B(n2699), .Y(n5864) );
  OAI21X1 U2658 ( .A(n4489), .B(n2697), .C(n5865), .Y(n8056) );
  NAND2X1 U2659 ( .A(arr[1298]), .B(n2699), .Y(n5865) );
  OAI21X1 U2660 ( .A(n4491), .B(n2698), .C(n5866), .Y(n8057) );
  NAND2X1 U2661 ( .A(arr[1299]), .B(n2699), .Y(n5866) );
  OAI21X1 U2662 ( .A(n4493), .B(n2698), .C(n5867), .Y(n8058) );
  NAND2X1 U2663 ( .A(arr[1300]), .B(n2699), .Y(n5867) );
  OAI21X1 U2664 ( .A(n4495), .B(n2697), .C(n5868), .Y(n8059) );
  NAND2X1 U2665 ( .A(arr[1301]), .B(n2699), .Y(n5868) );
  OAI21X1 U2666 ( .A(n4497), .B(n2698), .C(n5869), .Y(n8060) );
  NAND2X1 U2667 ( .A(arr[1302]), .B(n2699), .Y(n5869) );
  OAI21X1 U2668 ( .A(n4499), .B(n2698), .C(n5870), .Y(n8061) );
  NAND2X1 U2669 ( .A(arr[1303]), .B(n2699), .Y(n5870) );
  OAI21X1 U2670 ( .A(n4501), .B(n2697), .C(n5871), .Y(n8062) );
  NAND2X1 U2671 ( .A(arr[1304]), .B(n2699), .Y(n5871) );
  OAI21X1 U2672 ( .A(n4503), .B(n2697), .C(n5872), .Y(n8063) );
  NAND2X1 U2673 ( .A(arr[1305]), .B(n2699), .Y(n5872) );
  OAI21X1 U2674 ( .A(n4505), .B(n2697), .C(n5873), .Y(n8064) );
  NAND2X1 U2675 ( .A(arr[1306]), .B(n2699), .Y(n5873) );
  OAI21X1 U2676 ( .A(n4507), .B(n2697), .C(n5874), .Y(n8065) );
  NAND2X1 U2677 ( .A(arr[1307]), .B(n2699), .Y(n5874) );
  OAI21X1 U2678 ( .A(n4509), .B(n2697), .C(n5875), .Y(n8066) );
  NAND2X1 U2679 ( .A(arr[1308]), .B(n2699), .Y(n5875) );
  OAI21X1 U2680 ( .A(n4511), .B(n2697), .C(n5876), .Y(n8067) );
  NAND2X1 U2681 ( .A(arr[1309]), .B(n2699), .Y(n5876) );
  OAI21X1 U2682 ( .A(n4513), .B(n2699), .C(n5877), .Y(n8068) );
  NAND2X1 U2683 ( .A(arr[1310]), .B(n2699), .Y(n5877) );
  OAI21X1 U2684 ( .A(n4515), .B(n2697), .C(n5878), .Y(n8069) );
  NAND2X1 U2685 ( .A(arr[1311]), .B(n2699), .Y(n5878) );
  OAI21X1 U2686 ( .A(n4517), .B(n2698), .C(n5879), .Y(n8070) );
  NAND2X1 U2687 ( .A(arr[1312]), .B(n2699), .Y(n5879) );
  OAI21X1 U2688 ( .A(n4519), .B(n2697), .C(n5880), .Y(n8071) );
  NAND2X1 U2689 ( .A(arr[1313]), .B(n2698), .Y(n5880) );
  OAI21X1 U2690 ( .A(n4521), .B(n2698), .C(n5881), .Y(n8072) );
  NAND2X1 U2691 ( .A(arr[1314]), .B(n2699), .Y(n5881) );
  OAI21X1 U2692 ( .A(n4523), .B(n2697), .C(n5882), .Y(n8073) );
  NAND2X1 U2693 ( .A(arr[1315]), .B(n2698), .Y(n5882) );
  OAI21X1 U2694 ( .A(n4525), .B(n2697), .C(n5883), .Y(n8074) );
  NAND2X1 U2695 ( .A(arr[1316]), .B(n2699), .Y(n5883) );
  OAI21X1 U2696 ( .A(n4527), .B(n2697), .C(n5884), .Y(n8075) );
  NAND2X1 U2697 ( .A(arr[1317]), .B(n2698), .Y(n5884) );
  OAI21X1 U2698 ( .A(n4529), .B(n2697), .C(n5885), .Y(n8076) );
  NAND2X1 U2699 ( .A(arr[1318]), .B(n2698), .Y(n5885) );
  OAI21X1 U2700 ( .A(n4531), .B(n2697), .C(n5886), .Y(n8077) );
  NAND2X1 U2701 ( .A(arr[1319]), .B(n2699), .Y(n5886) );
  AND2X1 U2703 ( .A(n5887), .B(n5679), .Y(n4742) );
  NOR2X1 U2704 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .Y(n5679) );
  OAI21X1 U2705 ( .A(n4467), .B(n2696), .C(n5889), .Y(n8078) );
  NAND2X1 U2706 ( .A(arr[1320]), .B(n2695), .Y(n5889) );
  OAI21X1 U2707 ( .A(n4469), .B(n2694), .C(n5890), .Y(n8079) );
  NAND2X1 U2708 ( .A(arr[1321]), .B(n2695), .Y(n5890) );
  OAI21X1 U2709 ( .A(n4471), .B(n2694), .C(n5891), .Y(n8080) );
  NAND2X1 U2710 ( .A(arr[1322]), .B(n2695), .Y(n5891) );
  OAI21X1 U2711 ( .A(n4473), .B(n2694), .C(n5892), .Y(n8081) );
  NAND2X1 U2712 ( .A(arr[1323]), .B(n2695), .Y(n5892) );
  OAI21X1 U2713 ( .A(n4475), .B(n2694), .C(n5893), .Y(n8082) );
  NAND2X1 U2714 ( .A(arr[1324]), .B(n2695), .Y(n5893) );
  OAI21X1 U2715 ( .A(n4477), .B(n2694), .C(n5894), .Y(n8083) );
  NAND2X1 U2716 ( .A(arr[1325]), .B(n2696), .Y(n5894) );
  OAI21X1 U2717 ( .A(n4479), .B(n2694), .C(n5895), .Y(n8084) );
  NAND2X1 U2718 ( .A(arr[1326]), .B(n2696), .Y(n5895) );
  OAI21X1 U2719 ( .A(n4481), .B(n2695), .C(n5896), .Y(n8085) );
  NAND2X1 U2720 ( .A(arr[1327]), .B(n2695), .Y(n5896) );
  OAI21X1 U2721 ( .A(n4483), .B(n2694), .C(n5897), .Y(n8086) );
  NAND2X1 U2722 ( .A(arr[1328]), .B(n2695), .Y(n5897) );
  OAI21X1 U2723 ( .A(n4485), .B(n2695), .C(n5898), .Y(n8087) );
  NAND2X1 U2724 ( .A(arr[1329]), .B(n2696), .Y(n5898) );
  OAI21X1 U2725 ( .A(n4487), .B(n2695), .C(n5899), .Y(n8088) );
  NAND2X1 U2726 ( .A(arr[1330]), .B(n2696), .Y(n5899) );
  OAI21X1 U2727 ( .A(n4489), .B(n2694), .C(n5900), .Y(n8089) );
  NAND2X1 U2728 ( .A(arr[1331]), .B(n2696), .Y(n5900) );
  OAI21X1 U2729 ( .A(n4491), .B(n2695), .C(n5901), .Y(n8090) );
  NAND2X1 U2730 ( .A(arr[1332]), .B(n2696), .Y(n5901) );
  OAI21X1 U2731 ( .A(n4493), .B(n2695), .C(n5902), .Y(n8091) );
  NAND2X1 U2732 ( .A(arr[1333]), .B(n2696), .Y(n5902) );
  OAI21X1 U2733 ( .A(n4495), .B(n2694), .C(n5903), .Y(n8092) );
  NAND2X1 U2734 ( .A(arr[1334]), .B(n2696), .Y(n5903) );
  OAI21X1 U2735 ( .A(n4497), .B(n2695), .C(n5904), .Y(n8093) );
  NAND2X1 U2736 ( .A(arr[1335]), .B(n2696), .Y(n5904) );
  OAI21X1 U2737 ( .A(n4499), .B(n2695), .C(n5905), .Y(n8094) );
  NAND2X1 U2738 ( .A(arr[1336]), .B(n2696), .Y(n5905) );
  OAI21X1 U2739 ( .A(n4501), .B(n2694), .C(n5906), .Y(n8095) );
  NAND2X1 U2740 ( .A(arr[1337]), .B(n2696), .Y(n5906) );
  OAI21X1 U2741 ( .A(n4503), .B(n2694), .C(n5907), .Y(n8096) );
  NAND2X1 U2742 ( .A(arr[1338]), .B(n2696), .Y(n5907) );
  OAI21X1 U2743 ( .A(n4505), .B(n2694), .C(n5908), .Y(n8097) );
  NAND2X1 U2744 ( .A(arr[1339]), .B(n2696), .Y(n5908) );
  OAI21X1 U2745 ( .A(n4507), .B(n2694), .C(n5909), .Y(n8098) );
  NAND2X1 U2746 ( .A(arr[1340]), .B(n2696), .Y(n5909) );
  OAI21X1 U2747 ( .A(n4509), .B(n2694), .C(n5910), .Y(n8099) );
  NAND2X1 U2748 ( .A(arr[1341]), .B(n2696), .Y(n5910) );
  OAI21X1 U2749 ( .A(n4511), .B(n2694), .C(n5911), .Y(n8100) );
  NAND2X1 U2750 ( .A(arr[1342]), .B(n2696), .Y(n5911) );
  OAI21X1 U2751 ( .A(n4513), .B(n2696), .C(n5912), .Y(n8101) );
  NAND2X1 U2752 ( .A(arr[1343]), .B(n2696), .Y(n5912) );
  OAI21X1 U2753 ( .A(n4515), .B(n2694), .C(n5913), .Y(n8102) );
  NAND2X1 U2754 ( .A(arr[1344]), .B(n2696), .Y(n5913) );
  OAI21X1 U2755 ( .A(n4517), .B(n2695), .C(n5914), .Y(n8103) );
  NAND2X1 U2756 ( .A(arr[1345]), .B(n2696), .Y(n5914) );
  OAI21X1 U2757 ( .A(n4519), .B(n2694), .C(n5915), .Y(n8104) );
  NAND2X1 U2758 ( .A(arr[1346]), .B(n2695), .Y(n5915) );
  OAI21X1 U2759 ( .A(n4521), .B(n2695), .C(n5916), .Y(n8105) );
  NAND2X1 U2760 ( .A(arr[1347]), .B(n2696), .Y(n5916) );
  OAI21X1 U2761 ( .A(n4523), .B(n2694), .C(n5917), .Y(n8106) );
  NAND2X1 U2762 ( .A(arr[1348]), .B(n2695), .Y(n5917) );
  OAI21X1 U2763 ( .A(n4525), .B(n2694), .C(n5918), .Y(n8107) );
  NAND2X1 U2764 ( .A(arr[1349]), .B(n2696), .Y(n5918) );
  OAI21X1 U2765 ( .A(n4527), .B(n2694), .C(n5919), .Y(n8108) );
  NAND2X1 U2766 ( .A(arr[1350]), .B(n2695), .Y(n5919) );
  OAI21X1 U2767 ( .A(n4529), .B(n2694), .C(n5920), .Y(n8109) );
  NAND2X1 U2768 ( .A(arr[1351]), .B(n2695), .Y(n5920) );
  OAI21X1 U2769 ( .A(n4531), .B(n2694), .C(n5921), .Y(n8110) );
  NAND2X1 U2770 ( .A(arr[1352]), .B(n2696), .Y(n5921) );
  OAI21X1 U2772 ( .A(n4467), .B(n2693), .C(n5923), .Y(n8111) );
  NAND2X1 U2773 ( .A(arr[1353]), .B(n2692), .Y(n5923) );
  OAI21X1 U2774 ( .A(n4469), .B(n2691), .C(n5924), .Y(n8112) );
  NAND2X1 U2775 ( .A(arr[1354]), .B(n2692), .Y(n5924) );
  OAI21X1 U2776 ( .A(n4471), .B(n2691), .C(n5925), .Y(n8113) );
  NAND2X1 U2777 ( .A(arr[1355]), .B(n2692), .Y(n5925) );
  OAI21X1 U2778 ( .A(n4473), .B(n2691), .C(n5926), .Y(n8114) );
  NAND2X1 U2779 ( .A(arr[1356]), .B(n2692), .Y(n5926) );
  OAI21X1 U2780 ( .A(n4475), .B(n2691), .C(n5927), .Y(n8115) );
  NAND2X1 U2781 ( .A(arr[1357]), .B(n2692), .Y(n5927) );
  OAI21X1 U2782 ( .A(n4477), .B(n2691), .C(n5928), .Y(n8116) );
  NAND2X1 U2783 ( .A(arr[1358]), .B(n2693), .Y(n5928) );
  OAI21X1 U2784 ( .A(n4479), .B(n2691), .C(n5929), .Y(n8117) );
  NAND2X1 U2785 ( .A(arr[1359]), .B(n2693), .Y(n5929) );
  OAI21X1 U2786 ( .A(n4481), .B(n2692), .C(n5930), .Y(n8118) );
  NAND2X1 U2787 ( .A(arr[1360]), .B(n2692), .Y(n5930) );
  OAI21X1 U2788 ( .A(n4483), .B(n2691), .C(n5931), .Y(n8119) );
  NAND2X1 U2789 ( .A(arr[1361]), .B(n2692), .Y(n5931) );
  OAI21X1 U2790 ( .A(n4485), .B(n2692), .C(n5932), .Y(n8120) );
  NAND2X1 U2791 ( .A(arr[1362]), .B(n2693), .Y(n5932) );
  OAI21X1 U2792 ( .A(n4487), .B(n2692), .C(n5933), .Y(n8121) );
  NAND2X1 U2793 ( .A(arr[1363]), .B(n2693), .Y(n5933) );
  OAI21X1 U2794 ( .A(n4489), .B(n2691), .C(n5934), .Y(n8122) );
  NAND2X1 U2795 ( .A(arr[1364]), .B(n2693), .Y(n5934) );
  OAI21X1 U2796 ( .A(n4491), .B(n2692), .C(n5935), .Y(n8123) );
  NAND2X1 U2797 ( .A(arr[1365]), .B(n2693), .Y(n5935) );
  OAI21X1 U2798 ( .A(n4493), .B(n2692), .C(n5936), .Y(n8124) );
  NAND2X1 U2799 ( .A(arr[1366]), .B(n2693), .Y(n5936) );
  OAI21X1 U2800 ( .A(n4495), .B(n2691), .C(n5937), .Y(n8125) );
  NAND2X1 U2801 ( .A(arr[1367]), .B(n2693), .Y(n5937) );
  OAI21X1 U2802 ( .A(n4497), .B(n2692), .C(n5938), .Y(n8126) );
  NAND2X1 U2803 ( .A(arr[1368]), .B(n2693), .Y(n5938) );
  OAI21X1 U2804 ( .A(n4499), .B(n2692), .C(n5939), .Y(n8127) );
  NAND2X1 U2805 ( .A(arr[1369]), .B(n2693), .Y(n5939) );
  OAI21X1 U2806 ( .A(n4501), .B(n2691), .C(n5940), .Y(n8128) );
  NAND2X1 U2807 ( .A(arr[1370]), .B(n2693), .Y(n5940) );
  OAI21X1 U2808 ( .A(n4503), .B(n2691), .C(n5941), .Y(n8129) );
  NAND2X1 U2809 ( .A(arr[1371]), .B(n2693), .Y(n5941) );
  OAI21X1 U2810 ( .A(n4505), .B(n2691), .C(n5942), .Y(n8130) );
  NAND2X1 U2811 ( .A(arr[1372]), .B(n2693), .Y(n5942) );
  OAI21X1 U2812 ( .A(n4507), .B(n2691), .C(n5943), .Y(n8131) );
  NAND2X1 U2813 ( .A(arr[1373]), .B(n2693), .Y(n5943) );
  OAI21X1 U2814 ( .A(n4509), .B(n2691), .C(n5944), .Y(n8132) );
  NAND2X1 U2815 ( .A(arr[1374]), .B(n2693), .Y(n5944) );
  OAI21X1 U2816 ( .A(n4511), .B(n2691), .C(n5945), .Y(n8133) );
  NAND2X1 U2817 ( .A(arr[1375]), .B(n2693), .Y(n5945) );
  OAI21X1 U2818 ( .A(n4513), .B(n2693), .C(n5946), .Y(n8134) );
  NAND2X1 U2819 ( .A(arr[1376]), .B(n2693), .Y(n5946) );
  OAI21X1 U2820 ( .A(n4515), .B(n2691), .C(n5947), .Y(n8135) );
  NAND2X1 U2821 ( .A(arr[1377]), .B(n2693), .Y(n5947) );
  OAI21X1 U2822 ( .A(n4517), .B(n2692), .C(n5948), .Y(n8136) );
  NAND2X1 U2823 ( .A(arr[1378]), .B(n2693), .Y(n5948) );
  OAI21X1 U2824 ( .A(n4519), .B(n2691), .C(n5949), .Y(n8137) );
  NAND2X1 U2825 ( .A(arr[1379]), .B(n2692), .Y(n5949) );
  OAI21X1 U2826 ( .A(n4521), .B(n2692), .C(n5950), .Y(n8138) );
  NAND2X1 U2827 ( .A(arr[1380]), .B(n2693), .Y(n5950) );
  OAI21X1 U2828 ( .A(n4523), .B(n2691), .C(n5951), .Y(n8139) );
  NAND2X1 U2829 ( .A(arr[1381]), .B(n2692), .Y(n5951) );
  OAI21X1 U2830 ( .A(n4525), .B(n2691), .C(n5952), .Y(n8140) );
  NAND2X1 U2831 ( .A(arr[1382]), .B(n2693), .Y(n5952) );
  OAI21X1 U2832 ( .A(n4527), .B(n2691), .C(n5953), .Y(n8141) );
  NAND2X1 U2833 ( .A(arr[1383]), .B(n2692), .Y(n5953) );
  OAI21X1 U2834 ( .A(n4529), .B(n2691), .C(n5954), .Y(n8142) );
  NAND2X1 U2835 ( .A(arr[1384]), .B(n2692), .Y(n5954) );
  OAI21X1 U2836 ( .A(n4531), .B(n2691), .C(n5955), .Y(n8143) );
  NAND2X1 U2837 ( .A(arr[1385]), .B(n2693), .Y(n5955) );
  AND2X1 U2839 ( .A(n5956), .B(n5680), .Y(n4811) );
  OAI21X1 U2840 ( .A(n4467), .B(n2690), .C(n5958), .Y(n8144) );
  NAND2X1 U2841 ( .A(arr[1386]), .B(n2689), .Y(n5958) );
  OAI21X1 U2842 ( .A(n4469), .B(n2688), .C(n5959), .Y(n8145) );
  NAND2X1 U2843 ( .A(arr[1387]), .B(n2689), .Y(n5959) );
  OAI21X1 U2844 ( .A(n4471), .B(n2688), .C(n5960), .Y(n8146) );
  NAND2X1 U2845 ( .A(arr[1388]), .B(n2689), .Y(n5960) );
  OAI21X1 U2846 ( .A(n4473), .B(n2688), .C(n5961), .Y(n8147) );
  NAND2X1 U2847 ( .A(arr[1389]), .B(n2689), .Y(n5961) );
  OAI21X1 U2848 ( .A(n4475), .B(n2688), .C(n5962), .Y(n8148) );
  NAND2X1 U2849 ( .A(arr[1390]), .B(n2689), .Y(n5962) );
  OAI21X1 U2850 ( .A(n4477), .B(n2688), .C(n5963), .Y(n8149) );
  NAND2X1 U2851 ( .A(arr[1391]), .B(n2690), .Y(n5963) );
  OAI21X1 U2852 ( .A(n4479), .B(n2688), .C(n5964), .Y(n8150) );
  NAND2X1 U2853 ( .A(arr[1392]), .B(n2690), .Y(n5964) );
  OAI21X1 U2854 ( .A(n4481), .B(n2689), .C(n5965), .Y(n8151) );
  NAND2X1 U2855 ( .A(arr[1393]), .B(n2689), .Y(n5965) );
  OAI21X1 U2856 ( .A(n4483), .B(n2688), .C(n5966), .Y(n8152) );
  NAND2X1 U2857 ( .A(arr[1394]), .B(n2689), .Y(n5966) );
  OAI21X1 U2858 ( .A(n4485), .B(n2689), .C(n5967), .Y(n8153) );
  NAND2X1 U2859 ( .A(arr[1395]), .B(n2690), .Y(n5967) );
  OAI21X1 U2860 ( .A(n4487), .B(n2689), .C(n5968), .Y(n8154) );
  NAND2X1 U2861 ( .A(arr[1396]), .B(n2690), .Y(n5968) );
  OAI21X1 U2862 ( .A(n4489), .B(n2688), .C(n5969), .Y(n8155) );
  NAND2X1 U2863 ( .A(arr[1397]), .B(n2690), .Y(n5969) );
  OAI21X1 U2864 ( .A(n4491), .B(n2689), .C(n5970), .Y(n8156) );
  NAND2X1 U2865 ( .A(arr[1398]), .B(n2690), .Y(n5970) );
  OAI21X1 U2866 ( .A(n4493), .B(n2689), .C(n5971), .Y(n8157) );
  NAND2X1 U2867 ( .A(arr[1399]), .B(n2690), .Y(n5971) );
  OAI21X1 U2868 ( .A(n4495), .B(n2688), .C(n5972), .Y(n8158) );
  NAND2X1 U2869 ( .A(arr[1400]), .B(n2690), .Y(n5972) );
  OAI21X1 U2870 ( .A(n4497), .B(n2689), .C(n5973), .Y(n8159) );
  NAND2X1 U2871 ( .A(arr[1401]), .B(n2690), .Y(n5973) );
  OAI21X1 U2872 ( .A(n4499), .B(n2689), .C(n5974), .Y(n8160) );
  NAND2X1 U2873 ( .A(arr[1402]), .B(n2690), .Y(n5974) );
  OAI21X1 U2874 ( .A(n4501), .B(n2688), .C(n5975), .Y(n8161) );
  NAND2X1 U2875 ( .A(arr[1403]), .B(n2690), .Y(n5975) );
  OAI21X1 U2876 ( .A(n4503), .B(n2688), .C(n5976), .Y(n8162) );
  NAND2X1 U2877 ( .A(arr[1404]), .B(n2690), .Y(n5976) );
  OAI21X1 U2878 ( .A(n4505), .B(n2688), .C(n5977), .Y(n8163) );
  NAND2X1 U2879 ( .A(arr[1405]), .B(n2690), .Y(n5977) );
  OAI21X1 U2880 ( .A(n4507), .B(n2688), .C(n5978), .Y(n8164) );
  NAND2X1 U2881 ( .A(arr[1406]), .B(n2690), .Y(n5978) );
  OAI21X1 U2882 ( .A(n4509), .B(n2688), .C(n5979), .Y(n8165) );
  NAND2X1 U2883 ( .A(arr[1407]), .B(n2690), .Y(n5979) );
  OAI21X1 U2884 ( .A(n4511), .B(n2688), .C(n5980), .Y(n8166) );
  NAND2X1 U2885 ( .A(arr[1408]), .B(n2690), .Y(n5980) );
  OAI21X1 U2886 ( .A(n4513), .B(n2690), .C(n5981), .Y(n8167) );
  NAND2X1 U2887 ( .A(arr[1409]), .B(n2690), .Y(n5981) );
  OAI21X1 U2888 ( .A(n4515), .B(n2688), .C(n5982), .Y(n8168) );
  NAND2X1 U2889 ( .A(arr[1410]), .B(n2690), .Y(n5982) );
  OAI21X1 U2890 ( .A(n4517), .B(n2689), .C(n5983), .Y(n8169) );
  NAND2X1 U2891 ( .A(arr[1411]), .B(n2690), .Y(n5983) );
  OAI21X1 U2892 ( .A(n4519), .B(n2688), .C(n5984), .Y(n8170) );
  NAND2X1 U2893 ( .A(arr[1412]), .B(n2689), .Y(n5984) );
  OAI21X1 U2894 ( .A(n4521), .B(n2689), .C(n5985), .Y(n8171) );
  NAND2X1 U2895 ( .A(arr[1413]), .B(n2690), .Y(n5985) );
  OAI21X1 U2896 ( .A(n4523), .B(n2688), .C(n5986), .Y(n8172) );
  NAND2X1 U2897 ( .A(arr[1414]), .B(n2689), .Y(n5986) );
  OAI21X1 U2898 ( .A(n4525), .B(n2688), .C(n5987), .Y(n8173) );
  NAND2X1 U2899 ( .A(arr[1415]), .B(n2690), .Y(n5987) );
  OAI21X1 U2900 ( .A(n4527), .B(n2688), .C(n5988), .Y(n8174) );
  NAND2X1 U2901 ( .A(arr[1416]), .B(n2689), .Y(n5988) );
  OAI21X1 U2902 ( .A(n4529), .B(n2688), .C(n5989), .Y(n8175) );
  NAND2X1 U2903 ( .A(arr[1417]), .B(n2689), .Y(n5989) );
  OAI21X1 U2904 ( .A(n4531), .B(n2688), .C(n5990), .Y(n8176) );
  NAND2X1 U2905 ( .A(arr[1418]), .B(n2690), .Y(n5990) );
  OAI21X1 U2907 ( .A(n4467), .B(n2687), .C(n5992), .Y(n8177) );
  NAND2X1 U2908 ( .A(arr[1419]), .B(n2686), .Y(n5992) );
  OAI21X1 U2909 ( .A(n4469), .B(n2685), .C(n5993), .Y(n8178) );
  NAND2X1 U2910 ( .A(arr[1420]), .B(n2686), .Y(n5993) );
  OAI21X1 U2911 ( .A(n4471), .B(n2685), .C(n5994), .Y(n8179) );
  NAND2X1 U2912 ( .A(arr[1421]), .B(n2686), .Y(n5994) );
  OAI21X1 U2913 ( .A(n4473), .B(n2685), .C(n5995), .Y(n8180) );
  NAND2X1 U2914 ( .A(arr[1422]), .B(n2686), .Y(n5995) );
  OAI21X1 U2915 ( .A(n4475), .B(n2685), .C(n5996), .Y(n8181) );
  NAND2X1 U2916 ( .A(arr[1423]), .B(n2686), .Y(n5996) );
  OAI21X1 U2917 ( .A(n4477), .B(n2685), .C(n5997), .Y(n8182) );
  NAND2X1 U2918 ( .A(arr[1424]), .B(n2687), .Y(n5997) );
  OAI21X1 U2919 ( .A(n4479), .B(n2685), .C(n5998), .Y(n8183) );
  NAND2X1 U2920 ( .A(arr[1425]), .B(n2687), .Y(n5998) );
  OAI21X1 U2921 ( .A(n4481), .B(n2686), .C(n5999), .Y(n8184) );
  NAND2X1 U2922 ( .A(arr[1426]), .B(n2686), .Y(n5999) );
  OAI21X1 U2923 ( .A(n4483), .B(n2685), .C(n6000), .Y(n8185) );
  NAND2X1 U2924 ( .A(arr[1427]), .B(n2686), .Y(n6000) );
  OAI21X1 U2925 ( .A(n4485), .B(n2686), .C(n6001), .Y(n8186) );
  NAND2X1 U2926 ( .A(arr[1428]), .B(n2687), .Y(n6001) );
  OAI21X1 U2927 ( .A(n4487), .B(n2686), .C(n6002), .Y(n8187) );
  NAND2X1 U2928 ( .A(arr[1429]), .B(n2687), .Y(n6002) );
  OAI21X1 U2929 ( .A(n4489), .B(n2685), .C(n6003), .Y(n8188) );
  NAND2X1 U2930 ( .A(arr[1430]), .B(n2687), .Y(n6003) );
  OAI21X1 U2931 ( .A(n4491), .B(n2686), .C(n6004), .Y(n8189) );
  NAND2X1 U2932 ( .A(arr[1431]), .B(n2687), .Y(n6004) );
  OAI21X1 U2933 ( .A(n4493), .B(n2686), .C(n6005), .Y(n8190) );
  NAND2X1 U2934 ( .A(arr[1432]), .B(n2687), .Y(n6005) );
  OAI21X1 U2935 ( .A(n4495), .B(n2685), .C(n6006), .Y(n8191) );
  NAND2X1 U2936 ( .A(arr[1433]), .B(n2687), .Y(n6006) );
  OAI21X1 U2937 ( .A(n4497), .B(n2686), .C(n6007), .Y(n8192) );
  NAND2X1 U2938 ( .A(arr[1434]), .B(n2687), .Y(n6007) );
  OAI21X1 U2939 ( .A(n4499), .B(n2686), .C(n6008), .Y(n8193) );
  NAND2X1 U2940 ( .A(arr[1435]), .B(n2687), .Y(n6008) );
  OAI21X1 U2941 ( .A(n4501), .B(n2685), .C(n6009), .Y(n8194) );
  NAND2X1 U2942 ( .A(arr[1436]), .B(n2687), .Y(n6009) );
  OAI21X1 U2943 ( .A(n4503), .B(n2685), .C(n6010), .Y(n8195) );
  NAND2X1 U2944 ( .A(arr[1437]), .B(n2687), .Y(n6010) );
  OAI21X1 U2945 ( .A(n4505), .B(n2685), .C(n6011), .Y(n8196) );
  NAND2X1 U2946 ( .A(arr[1438]), .B(n2687), .Y(n6011) );
  OAI21X1 U2947 ( .A(n4507), .B(n2685), .C(n6012), .Y(n8197) );
  NAND2X1 U2948 ( .A(arr[1439]), .B(n2687), .Y(n6012) );
  OAI21X1 U2949 ( .A(n4509), .B(n2685), .C(n6013), .Y(n8198) );
  NAND2X1 U2950 ( .A(arr[1440]), .B(n2687), .Y(n6013) );
  OAI21X1 U2951 ( .A(n4511), .B(n2685), .C(n6014), .Y(n8199) );
  NAND2X1 U2952 ( .A(arr[1441]), .B(n2687), .Y(n6014) );
  OAI21X1 U2953 ( .A(n4513), .B(n2687), .C(n6015), .Y(n8200) );
  NAND2X1 U2954 ( .A(arr[1442]), .B(n2687), .Y(n6015) );
  OAI21X1 U2955 ( .A(n4515), .B(n2685), .C(n6016), .Y(n8201) );
  NAND2X1 U2956 ( .A(arr[1443]), .B(n2687), .Y(n6016) );
  OAI21X1 U2957 ( .A(n4517), .B(n2686), .C(n6017), .Y(n8202) );
  NAND2X1 U2958 ( .A(arr[1444]), .B(n2687), .Y(n6017) );
  OAI21X1 U2959 ( .A(n4519), .B(n2685), .C(n6018), .Y(n8203) );
  NAND2X1 U2960 ( .A(arr[1445]), .B(n2686), .Y(n6018) );
  OAI21X1 U2961 ( .A(n4521), .B(n2686), .C(n6019), .Y(n8204) );
  NAND2X1 U2962 ( .A(arr[1446]), .B(n2687), .Y(n6019) );
  OAI21X1 U2963 ( .A(n4523), .B(n2685), .C(n6020), .Y(n8205) );
  NAND2X1 U2964 ( .A(arr[1447]), .B(n2686), .Y(n6020) );
  OAI21X1 U2965 ( .A(n4525), .B(n2685), .C(n6021), .Y(n8206) );
  NAND2X1 U2966 ( .A(arr[1448]), .B(n2687), .Y(n6021) );
  OAI21X1 U2967 ( .A(n4527), .B(n2685), .C(n6022), .Y(n8207) );
  NAND2X1 U2968 ( .A(arr[1449]), .B(n2686), .Y(n6022) );
  OAI21X1 U2969 ( .A(n4529), .B(n2685), .C(n6023), .Y(n8208) );
  NAND2X1 U2970 ( .A(arr[1450]), .B(n2686), .Y(n6023) );
  OAI21X1 U2971 ( .A(n4531), .B(n2685), .C(n6024), .Y(n8209) );
  NAND2X1 U2972 ( .A(arr[1451]), .B(n2687), .Y(n6024) );
  AND2X1 U2974 ( .A(n5956), .B(n5749), .Y(n4880) );
  OAI21X1 U2975 ( .A(n4467), .B(n2684), .C(n6026), .Y(n8210) );
  NAND2X1 U2976 ( .A(arr[1452]), .B(n2683), .Y(n6026) );
  OAI21X1 U2977 ( .A(n4469), .B(n2682), .C(n6027), .Y(n8211) );
  NAND2X1 U2978 ( .A(arr[1453]), .B(n2683), .Y(n6027) );
  OAI21X1 U2979 ( .A(n4471), .B(n2682), .C(n6028), .Y(n8212) );
  NAND2X1 U2980 ( .A(arr[1454]), .B(n2683), .Y(n6028) );
  OAI21X1 U2981 ( .A(n4473), .B(n2682), .C(n6029), .Y(n8213) );
  NAND2X1 U2982 ( .A(arr[1455]), .B(n2683), .Y(n6029) );
  OAI21X1 U2983 ( .A(n4475), .B(n2682), .C(n6030), .Y(n8214) );
  NAND2X1 U2984 ( .A(arr[1456]), .B(n2683), .Y(n6030) );
  OAI21X1 U2985 ( .A(n4477), .B(n2682), .C(n6031), .Y(n8215) );
  NAND2X1 U2986 ( .A(arr[1457]), .B(n2684), .Y(n6031) );
  OAI21X1 U2987 ( .A(n4479), .B(n2682), .C(n6032), .Y(n8216) );
  NAND2X1 U2988 ( .A(arr[1458]), .B(n2684), .Y(n6032) );
  OAI21X1 U2989 ( .A(n4481), .B(n2683), .C(n6033), .Y(n8217) );
  NAND2X1 U2990 ( .A(arr[1459]), .B(n2683), .Y(n6033) );
  OAI21X1 U2991 ( .A(n4483), .B(n2682), .C(n6034), .Y(n8218) );
  NAND2X1 U2992 ( .A(arr[1460]), .B(n2683), .Y(n6034) );
  OAI21X1 U2993 ( .A(n4485), .B(n2683), .C(n6035), .Y(n8219) );
  NAND2X1 U2994 ( .A(arr[1461]), .B(n2684), .Y(n6035) );
  OAI21X1 U2995 ( .A(n4487), .B(n2683), .C(n6036), .Y(n8220) );
  NAND2X1 U2996 ( .A(arr[1462]), .B(n2684), .Y(n6036) );
  OAI21X1 U2997 ( .A(n4489), .B(n2682), .C(n6037), .Y(n8221) );
  NAND2X1 U2998 ( .A(arr[1463]), .B(n2684), .Y(n6037) );
  OAI21X1 U2999 ( .A(n4491), .B(n2683), .C(n6038), .Y(n8222) );
  NAND2X1 U3000 ( .A(arr[1464]), .B(n2684), .Y(n6038) );
  OAI21X1 U3001 ( .A(n4493), .B(n2683), .C(n6039), .Y(n8223) );
  NAND2X1 U3002 ( .A(arr[1465]), .B(n2684), .Y(n6039) );
  OAI21X1 U3003 ( .A(n4495), .B(n2682), .C(n6040), .Y(n8224) );
  NAND2X1 U3004 ( .A(arr[1466]), .B(n2684), .Y(n6040) );
  OAI21X1 U3005 ( .A(n4497), .B(n2683), .C(n6041), .Y(n8225) );
  NAND2X1 U3006 ( .A(arr[1467]), .B(n2684), .Y(n6041) );
  OAI21X1 U3007 ( .A(n4499), .B(n2683), .C(n6042), .Y(n8226) );
  NAND2X1 U3008 ( .A(arr[1468]), .B(n2684), .Y(n6042) );
  OAI21X1 U3009 ( .A(n4501), .B(n2682), .C(n6043), .Y(n8227) );
  NAND2X1 U3010 ( .A(arr[1469]), .B(n2684), .Y(n6043) );
  OAI21X1 U3011 ( .A(n4503), .B(n2682), .C(n6044), .Y(n8228) );
  NAND2X1 U3012 ( .A(arr[1470]), .B(n2684), .Y(n6044) );
  OAI21X1 U3013 ( .A(n4505), .B(n2682), .C(n6045), .Y(n8229) );
  NAND2X1 U3014 ( .A(arr[1471]), .B(n2684), .Y(n6045) );
  OAI21X1 U3015 ( .A(n4507), .B(n2682), .C(n6046), .Y(n8230) );
  NAND2X1 U3016 ( .A(arr[1472]), .B(n2684), .Y(n6046) );
  OAI21X1 U3017 ( .A(n4509), .B(n2682), .C(n6047), .Y(n8231) );
  NAND2X1 U3018 ( .A(arr[1473]), .B(n2684), .Y(n6047) );
  OAI21X1 U3019 ( .A(n4511), .B(n2682), .C(n6048), .Y(n8232) );
  NAND2X1 U3020 ( .A(arr[1474]), .B(n2684), .Y(n6048) );
  OAI21X1 U3021 ( .A(n4513), .B(n2684), .C(n6049), .Y(n8233) );
  NAND2X1 U3022 ( .A(arr[1475]), .B(n2684), .Y(n6049) );
  OAI21X1 U3023 ( .A(n4515), .B(n2682), .C(n6050), .Y(n8234) );
  NAND2X1 U3024 ( .A(arr[1476]), .B(n2684), .Y(n6050) );
  OAI21X1 U3025 ( .A(n4517), .B(n2683), .C(n6051), .Y(n8235) );
  NAND2X1 U3026 ( .A(arr[1477]), .B(n2684), .Y(n6051) );
  OAI21X1 U3027 ( .A(n4519), .B(n2682), .C(n6052), .Y(n8236) );
  NAND2X1 U3028 ( .A(arr[1478]), .B(n2683), .Y(n6052) );
  OAI21X1 U3029 ( .A(n4521), .B(n2683), .C(n6053), .Y(n8237) );
  NAND2X1 U3030 ( .A(arr[1479]), .B(n2684), .Y(n6053) );
  OAI21X1 U3031 ( .A(n4523), .B(n2682), .C(n6054), .Y(n8238) );
  NAND2X1 U3032 ( .A(arr[1480]), .B(n2683), .Y(n6054) );
  OAI21X1 U3033 ( .A(n4525), .B(n2682), .C(n6055), .Y(n8239) );
  NAND2X1 U3034 ( .A(arr[1481]), .B(n2684), .Y(n6055) );
  OAI21X1 U3035 ( .A(n4527), .B(n2682), .C(n6056), .Y(n8240) );
  NAND2X1 U3036 ( .A(arr[1482]), .B(n2683), .Y(n6056) );
  OAI21X1 U3037 ( .A(n4529), .B(n2682), .C(n6057), .Y(n8241) );
  NAND2X1 U3038 ( .A(arr[1483]), .B(n2683), .Y(n6057) );
  OAI21X1 U3039 ( .A(n4531), .B(n2682), .C(n6058), .Y(n8242) );
  NAND2X1 U3040 ( .A(arr[1484]), .B(n2684), .Y(n6058) );
  OAI21X1 U3042 ( .A(n4467), .B(n2681), .C(n6060), .Y(n8243) );
  NAND2X1 U3043 ( .A(arr[1485]), .B(n2680), .Y(n6060) );
  OAI21X1 U3044 ( .A(n4469), .B(n2679), .C(n6061), .Y(n8244) );
  NAND2X1 U3045 ( .A(arr[1486]), .B(n2680), .Y(n6061) );
  OAI21X1 U3046 ( .A(n4471), .B(n2679), .C(n6062), .Y(n8245) );
  NAND2X1 U3047 ( .A(arr[1487]), .B(n2680), .Y(n6062) );
  OAI21X1 U3048 ( .A(n4473), .B(n2679), .C(n6063), .Y(n8246) );
  NAND2X1 U3049 ( .A(arr[1488]), .B(n2680), .Y(n6063) );
  OAI21X1 U3050 ( .A(n4475), .B(n2679), .C(n6064), .Y(n8247) );
  NAND2X1 U3051 ( .A(arr[1489]), .B(n2680), .Y(n6064) );
  OAI21X1 U3052 ( .A(n4477), .B(n2679), .C(n6065), .Y(n8248) );
  NAND2X1 U3053 ( .A(arr[1490]), .B(n2681), .Y(n6065) );
  OAI21X1 U3054 ( .A(n4479), .B(n2679), .C(n6066), .Y(n8249) );
  NAND2X1 U3055 ( .A(arr[1491]), .B(n2681), .Y(n6066) );
  OAI21X1 U3056 ( .A(n4481), .B(n2680), .C(n6067), .Y(n8250) );
  NAND2X1 U3057 ( .A(arr[1492]), .B(n2680), .Y(n6067) );
  OAI21X1 U3058 ( .A(n4483), .B(n2679), .C(n6068), .Y(n8251) );
  NAND2X1 U3059 ( .A(arr[1493]), .B(n2680), .Y(n6068) );
  OAI21X1 U3060 ( .A(n4485), .B(n2680), .C(n6069), .Y(n8252) );
  NAND2X1 U3061 ( .A(arr[1494]), .B(n2681), .Y(n6069) );
  OAI21X1 U3062 ( .A(n4487), .B(n2680), .C(n6070), .Y(n8253) );
  NAND2X1 U3063 ( .A(arr[1495]), .B(n2681), .Y(n6070) );
  OAI21X1 U3064 ( .A(n4489), .B(n2679), .C(n6071), .Y(n8254) );
  NAND2X1 U3065 ( .A(arr[1496]), .B(n2681), .Y(n6071) );
  OAI21X1 U3066 ( .A(n4491), .B(n2680), .C(n6072), .Y(n8255) );
  NAND2X1 U3067 ( .A(arr[1497]), .B(n2681), .Y(n6072) );
  OAI21X1 U3068 ( .A(n4493), .B(n2680), .C(n6073), .Y(n8256) );
  NAND2X1 U3069 ( .A(arr[1498]), .B(n2681), .Y(n6073) );
  OAI21X1 U3070 ( .A(n4495), .B(n2679), .C(n6074), .Y(n8257) );
  NAND2X1 U3071 ( .A(arr[1499]), .B(n2681), .Y(n6074) );
  OAI21X1 U3072 ( .A(n4497), .B(n2680), .C(n6075), .Y(n8258) );
  NAND2X1 U3073 ( .A(arr[1500]), .B(n2681), .Y(n6075) );
  OAI21X1 U3074 ( .A(n4499), .B(n2680), .C(n6076), .Y(n8259) );
  NAND2X1 U3075 ( .A(arr[1501]), .B(n2681), .Y(n6076) );
  OAI21X1 U3076 ( .A(n4501), .B(n2679), .C(n6077), .Y(n8260) );
  NAND2X1 U3077 ( .A(arr[1502]), .B(n2681), .Y(n6077) );
  OAI21X1 U3078 ( .A(n4503), .B(n2679), .C(n6078), .Y(n8261) );
  NAND2X1 U3079 ( .A(arr[1503]), .B(n2681), .Y(n6078) );
  OAI21X1 U3080 ( .A(n4505), .B(n2679), .C(n6079), .Y(n8262) );
  NAND2X1 U3081 ( .A(arr[1504]), .B(n2681), .Y(n6079) );
  OAI21X1 U3082 ( .A(n4507), .B(n2679), .C(n6080), .Y(n8263) );
  NAND2X1 U3083 ( .A(arr[1505]), .B(n2681), .Y(n6080) );
  OAI21X1 U3084 ( .A(n4509), .B(n2679), .C(n6081), .Y(n8264) );
  NAND2X1 U3085 ( .A(arr[1506]), .B(n2681), .Y(n6081) );
  OAI21X1 U3086 ( .A(n4511), .B(n2679), .C(n6082), .Y(n8265) );
  NAND2X1 U3087 ( .A(arr[1507]), .B(n2681), .Y(n6082) );
  OAI21X1 U3088 ( .A(n4513), .B(n2681), .C(n6083), .Y(n8266) );
  NAND2X1 U3089 ( .A(arr[1508]), .B(n2681), .Y(n6083) );
  OAI21X1 U3090 ( .A(n4515), .B(n2679), .C(n6084), .Y(n8267) );
  NAND2X1 U3091 ( .A(arr[1509]), .B(n2681), .Y(n6084) );
  OAI21X1 U3092 ( .A(n4517), .B(n2680), .C(n6085), .Y(n8268) );
  NAND2X1 U3093 ( .A(arr[1510]), .B(n2681), .Y(n6085) );
  OAI21X1 U3094 ( .A(n4519), .B(n2679), .C(n6086), .Y(n8269) );
  NAND2X1 U3095 ( .A(arr[1511]), .B(n2680), .Y(n6086) );
  OAI21X1 U3096 ( .A(n4521), .B(n2680), .C(n6087), .Y(n8270) );
  NAND2X1 U3097 ( .A(arr[1512]), .B(n2681), .Y(n6087) );
  OAI21X1 U3098 ( .A(n4523), .B(n2679), .C(n6088), .Y(n8271) );
  NAND2X1 U3099 ( .A(arr[1513]), .B(n2680), .Y(n6088) );
  OAI21X1 U3100 ( .A(n4525), .B(n2679), .C(n6089), .Y(n8272) );
  NAND2X1 U3101 ( .A(arr[1514]), .B(n2681), .Y(n6089) );
  OAI21X1 U3102 ( .A(n4527), .B(n2679), .C(n6090), .Y(n8273) );
  NAND2X1 U3103 ( .A(arr[1515]), .B(n2680), .Y(n6090) );
  OAI21X1 U3104 ( .A(n4529), .B(n2679), .C(n6091), .Y(n8274) );
  NAND2X1 U3105 ( .A(arr[1516]), .B(n2680), .Y(n6091) );
  OAI21X1 U3106 ( .A(n4531), .B(n2679), .C(n6092), .Y(n8275) );
  NAND2X1 U3107 ( .A(arr[1517]), .B(n2681), .Y(n6092) );
  AND2X1 U3109 ( .A(n5956), .B(n5818), .Y(n4949) );
  OAI21X1 U3110 ( .A(n4467), .B(n2678), .C(n6094), .Y(n8276) );
  NAND2X1 U3111 ( .A(arr[1518]), .B(n2677), .Y(n6094) );
  OAI21X1 U3112 ( .A(n4469), .B(n2676), .C(n6095), .Y(n8277) );
  NAND2X1 U3113 ( .A(arr[1519]), .B(n2677), .Y(n6095) );
  OAI21X1 U3114 ( .A(n4471), .B(n2676), .C(n6096), .Y(n8278) );
  NAND2X1 U3115 ( .A(arr[1520]), .B(n2677), .Y(n6096) );
  OAI21X1 U3116 ( .A(n4473), .B(n2676), .C(n6097), .Y(n8279) );
  NAND2X1 U3117 ( .A(arr[1521]), .B(n2677), .Y(n6097) );
  OAI21X1 U3118 ( .A(n4475), .B(n2676), .C(n6098), .Y(n8280) );
  NAND2X1 U3119 ( .A(arr[1522]), .B(n2677), .Y(n6098) );
  OAI21X1 U3120 ( .A(n4477), .B(n2676), .C(n6099), .Y(n8281) );
  NAND2X1 U3121 ( .A(arr[1523]), .B(n2678), .Y(n6099) );
  OAI21X1 U3122 ( .A(n4479), .B(n2676), .C(n6100), .Y(n8282) );
  NAND2X1 U3123 ( .A(arr[1524]), .B(n2678), .Y(n6100) );
  OAI21X1 U3124 ( .A(n4481), .B(n2677), .C(n6101), .Y(n8283) );
  NAND2X1 U3125 ( .A(arr[1525]), .B(n2677), .Y(n6101) );
  OAI21X1 U3126 ( .A(n4483), .B(n2676), .C(n6102), .Y(n8284) );
  NAND2X1 U3127 ( .A(arr[1526]), .B(n2677), .Y(n6102) );
  OAI21X1 U3128 ( .A(n4485), .B(n2677), .C(n6103), .Y(n8285) );
  NAND2X1 U3129 ( .A(arr[1527]), .B(n2678), .Y(n6103) );
  OAI21X1 U3130 ( .A(n4487), .B(n2677), .C(n6104), .Y(n8286) );
  NAND2X1 U3131 ( .A(arr[1528]), .B(n2678), .Y(n6104) );
  OAI21X1 U3132 ( .A(n4489), .B(n2676), .C(n6105), .Y(n8287) );
  NAND2X1 U3133 ( .A(arr[1529]), .B(n2678), .Y(n6105) );
  OAI21X1 U3134 ( .A(n4491), .B(n2677), .C(n6106), .Y(n8288) );
  NAND2X1 U3135 ( .A(arr[1530]), .B(n2678), .Y(n6106) );
  OAI21X1 U3136 ( .A(n4493), .B(n2677), .C(n6107), .Y(n8289) );
  NAND2X1 U3137 ( .A(arr[1531]), .B(n2678), .Y(n6107) );
  OAI21X1 U3138 ( .A(n4495), .B(n2676), .C(n6108), .Y(n8290) );
  NAND2X1 U3139 ( .A(arr[1532]), .B(n2678), .Y(n6108) );
  OAI21X1 U3140 ( .A(n4497), .B(n2677), .C(n6109), .Y(n8291) );
  NAND2X1 U3141 ( .A(arr[1533]), .B(n2678), .Y(n6109) );
  OAI21X1 U3142 ( .A(n4499), .B(n2677), .C(n6110), .Y(n8292) );
  NAND2X1 U3143 ( .A(arr[1534]), .B(n2678), .Y(n6110) );
  OAI21X1 U3144 ( .A(n4501), .B(n2676), .C(n6111), .Y(n8293) );
  NAND2X1 U3145 ( .A(arr[1535]), .B(n2678), .Y(n6111) );
  OAI21X1 U3146 ( .A(n4503), .B(n2676), .C(n6112), .Y(n8294) );
  NAND2X1 U3147 ( .A(arr[1536]), .B(n2678), .Y(n6112) );
  OAI21X1 U3148 ( .A(n4505), .B(n2676), .C(n6113), .Y(n8295) );
  NAND2X1 U3149 ( .A(arr[1537]), .B(n2678), .Y(n6113) );
  OAI21X1 U3150 ( .A(n4507), .B(n2676), .C(n6114), .Y(n8296) );
  NAND2X1 U3151 ( .A(arr[1538]), .B(n2678), .Y(n6114) );
  OAI21X1 U3152 ( .A(n4509), .B(n2676), .C(n6115), .Y(n8297) );
  NAND2X1 U3153 ( .A(arr[1539]), .B(n2678), .Y(n6115) );
  OAI21X1 U3154 ( .A(n4511), .B(n2676), .C(n6116), .Y(n8298) );
  NAND2X1 U3155 ( .A(arr[1540]), .B(n2678), .Y(n6116) );
  OAI21X1 U3156 ( .A(n4513), .B(n2678), .C(n6117), .Y(n8299) );
  NAND2X1 U3157 ( .A(arr[1541]), .B(n2678), .Y(n6117) );
  OAI21X1 U3158 ( .A(n4515), .B(n2676), .C(n6118), .Y(n8300) );
  NAND2X1 U3159 ( .A(arr[1542]), .B(n2678), .Y(n6118) );
  OAI21X1 U3160 ( .A(n4517), .B(n2677), .C(n6119), .Y(n8301) );
  NAND2X1 U3161 ( .A(arr[1543]), .B(n2678), .Y(n6119) );
  OAI21X1 U3162 ( .A(n4519), .B(n2676), .C(n6120), .Y(n8302) );
  NAND2X1 U3163 ( .A(arr[1544]), .B(n2677), .Y(n6120) );
  OAI21X1 U3164 ( .A(n4521), .B(n2677), .C(n6121), .Y(n8303) );
  NAND2X1 U3165 ( .A(arr[1545]), .B(n2678), .Y(n6121) );
  OAI21X1 U3166 ( .A(n4523), .B(n2676), .C(n6122), .Y(n8304) );
  NAND2X1 U3167 ( .A(arr[1546]), .B(n2677), .Y(n6122) );
  OAI21X1 U3168 ( .A(n4525), .B(n2676), .C(n6123), .Y(n8305) );
  NAND2X1 U3169 ( .A(arr[1547]), .B(n2678), .Y(n6123) );
  OAI21X1 U3170 ( .A(n4527), .B(n2676), .C(n6124), .Y(n8306) );
  NAND2X1 U3171 ( .A(arr[1548]), .B(n2677), .Y(n6124) );
  OAI21X1 U3172 ( .A(n4529), .B(n2676), .C(n6125), .Y(n8307) );
  NAND2X1 U3173 ( .A(arr[1549]), .B(n2677), .Y(n6125) );
  OAI21X1 U3174 ( .A(n4531), .B(n2676), .C(n6126), .Y(n8308) );
  NAND2X1 U3175 ( .A(arr[1550]), .B(n2678), .Y(n6126) );
  OAI21X1 U3177 ( .A(n4467), .B(n2675), .C(n6128), .Y(n8309) );
  NAND2X1 U3178 ( .A(arr[1551]), .B(n2674), .Y(n6128) );
  OAI21X1 U3179 ( .A(n4469), .B(n2673), .C(n6129), .Y(n8310) );
  NAND2X1 U3180 ( .A(arr[1552]), .B(n2674), .Y(n6129) );
  OAI21X1 U3181 ( .A(n4471), .B(n2673), .C(n6130), .Y(n8311) );
  NAND2X1 U3182 ( .A(arr[1553]), .B(n2674), .Y(n6130) );
  OAI21X1 U3183 ( .A(n4473), .B(n2673), .C(n6131), .Y(n8312) );
  NAND2X1 U3184 ( .A(arr[1554]), .B(n2674), .Y(n6131) );
  OAI21X1 U3185 ( .A(n4475), .B(n2673), .C(n6132), .Y(n8313) );
  NAND2X1 U3186 ( .A(arr[1555]), .B(n2674), .Y(n6132) );
  OAI21X1 U3187 ( .A(n4477), .B(n2673), .C(n6133), .Y(n8314) );
  NAND2X1 U3188 ( .A(arr[1556]), .B(n2675), .Y(n6133) );
  OAI21X1 U3189 ( .A(n4479), .B(n2673), .C(n6134), .Y(n8315) );
  NAND2X1 U3190 ( .A(arr[1557]), .B(n2675), .Y(n6134) );
  OAI21X1 U3191 ( .A(n4481), .B(n2674), .C(n6135), .Y(n8316) );
  NAND2X1 U3192 ( .A(arr[1558]), .B(n2674), .Y(n6135) );
  OAI21X1 U3193 ( .A(n4483), .B(n2673), .C(n6136), .Y(n8317) );
  NAND2X1 U3194 ( .A(arr[1559]), .B(n2674), .Y(n6136) );
  OAI21X1 U3195 ( .A(n4485), .B(n2674), .C(n6137), .Y(n8318) );
  NAND2X1 U3196 ( .A(arr[1560]), .B(n2675), .Y(n6137) );
  OAI21X1 U3197 ( .A(n4487), .B(n2674), .C(n6138), .Y(n8319) );
  NAND2X1 U3198 ( .A(arr[1561]), .B(n2675), .Y(n6138) );
  OAI21X1 U3199 ( .A(n4489), .B(n2673), .C(n6139), .Y(n8320) );
  NAND2X1 U3200 ( .A(arr[1562]), .B(n2675), .Y(n6139) );
  OAI21X1 U3201 ( .A(n4491), .B(n2674), .C(n6140), .Y(n8321) );
  NAND2X1 U3202 ( .A(arr[1563]), .B(n2675), .Y(n6140) );
  OAI21X1 U3203 ( .A(n4493), .B(n2674), .C(n6141), .Y(n8322) );
  NAND2X1 U3204 ( .A(arr[1564]), .B(n2675), .Y(n6141) );
  OAI21X1 U3205 ( .A(n4495), .B(n2673), .C(n6142), .Y(n8323) );
  NAND2X1 U3206 ( .A(arr[1565]), .B(n2675), .Y(n6142) );
  OAI21X1 U3207 ( .A(n4497), .B(n2674), .C(n6143), .Y(n8324) );
  NAND2X1 U3208 ( .A(arr[1566]), .B(n2675), .Y(n6143) );
  OAI21X1 U3209 ( .A(n4499), .B(n2674), .C(n6144), .Y(n8325) );
  NAND2X1 U3210 ( .A(arr[1567]), .B(n2675), .Y(n6144) );
  OAI21X1 U3211 ( .A(n4501), .B(n2673), .C(n6145), .Y(n8326) );
  NAND2X1 U3212 ( .A(arr[1568]), .B(n2675), .Y(n6145) );
  OAI21X1 U3213 ( .A(n4503), .B(n2673), .C(n6146), .Y(n8327) );
  NAND2X1 U3214 ( .A(arr[1569]), .B(n2675), .Y(n6146) );
  OAI21X1 U3215 ( .A(n4505), .B(n2673), .C(n6147), .Y(n8328) );
  NAND2X1 U3216 ( .A(arr[1570]), .B(n2675), .Y(n6147) );
  OAI21X1 U3217 ( .A(n4507), .B(n2673), .C(n6148), .Y(n8329) );
  NAND2X1 U3218 ( .A(arr[1571]), .B(n2675), .Y(n6148) );
  OAI21X1 U3219 ( .A(n4509), .B(n2673), .C(n6149), .Y(n8330) );
  NAND2X1 U3220 ( .A(arr[1572]), .B(n2675), .Y(n6149) );
  OAI21X1 U3221 ( .A(n4511), .B(n2673), .C(n6150), .Y(n8331) );
  NAND2X1 U3222 ( .A(arr[1573]), .B(n2675), .Y(n6150) );
  OAI21X1 U3223 ( .A(n4513), .B(n2675), .C(n6151), .Y(n8332) );
  NAND2X1 U3224 ( .A(arr[1574]), .B(n2675), .Y(n6151) );
  OAI21X1 U3225 ( .A(n4515), .B(n2673), .C(n6152), .Y(n8333) );
  NAND2X1 U3226 ( .A(arr[1575]), .B(n2675), .Y(n6152) );
  OAI21X1 U3227 ( .A(n4517), .B(n2674), .C(n6153), .Y(n8334) );
  NAND2X1 U3228 ( .A(arr[1576]), .B(n2675), .Y(n6153) );
  OAI21X1 U3229 ( .A(n4519), .B(n2673), .C(n6154), .Y(n8335) );
  NAND2X1 U3230 ( .A(arr[1577]), .B(n2674), .Y(n6154) );
  OAI21X1 U3231 ( .A(n4521), .B(n2674), .C(n6155), .Y(n8336) );
  NAND2X1 U3232 ( .A(arr[1578]), .B(n2675), .Y(n6155) );
  OAI21X1 U3233 ( .A(n4523), .B(n2673), .C(n6156), .Y(n8337) );
  NAND2X1 U3234 ( .A(arr[1579]), .B(n2674), .Y(n6156) );
  OAI21X1 U3235 ( .A(n4525), .B(n2673), .C(n6157), .Y(n8338) );
  NAND2X1 U3236 ( .A(arr[1580]), .B(n2675), .Y(n6157) );
  OAI21X1 U3237 ( .A(n4527), .B(n2673), .C(n6158), .Y(n8339) );
  NAND2X1 U3238 ( .A(arr[1581]), .B(n2674), .Y(n6158) );
  OAI21X1 U3239 ( .A(n4529), .B(n2673), .C(n6159), .Y(n8340) );
  NAND2X1 U3240 ( .A(arr[1582]), .B(n2674), .Y(n6159) );
  OAI21X1 U3241 ( .A(n4531), .B(n2673), .C(n6160), .Y(n8341) );
  NAND2X1 U3242 ( .A(arr[1583]), .B(n2675), .Y(n6160) );
  AND2X1 U3244 ( .A(n5956), .B(n5887), .Y(n5018) );
  NOR2X1 U3245 ( .A(n6161), .B(wr_ptr[4]), .Y(n5956) );
  OAI21X1 U3246 ( .A(n4467), .B(n2672), .C(n6163), .Y(n8342) );
  NAND2X1 U3247 ( .A(arr[1584]), .B(n2671), .Y(n6163) );
  OAI21X1 U3248 ( .A(n4469), .B(n2670), .C(n6164), .Y(n8343) );
  NAND2X1 U3249 ( .A(arr[1585]), .B(n2671), .Y(n6164) );
  OAI21X1 U3250 ( .A(n4471), .B(n2670), .C(n6165), .Y(n8344) );
  NAND2X1 U3251 ( .A(arr[1586]), .B(n2671), .Y(n6165) );
  OAI21X1 U3252 ( .A(n4473), .B(n2670), .C(n6166), .Y(n8345) );
  NAND2X1 U3253 ( .A(arr[1587]), .B(n2671), .Y(n6166) );
  OAI21X1 U3254 ( .A(n4475), .B(n2670), .C(n6167), .Y(n8346) );
  NAND2X1 U3255 ( .A(arr[1588]), .B(n2671), .Y(n6167) );
  OAI21X1 U3256 ( .A(n4477), .B(n2670), .C(n6168), .Y(n8347) );
  NAND2X1 U3257 ( .A(arr[1589]), .B(n2672), .Y(n6168) );
  OAI21X1 U3258 ( .A(n4479), .B(n2670), .C(n6169), .Y(n8348) );
  NAND2X1 U3259 ( .A(arr[1590]), .B(n2672), .Y(n6169) );
  OAI21X1 U3260 ( .A(n4481), .B(n2671), .C(n6170), .Y(n8349) );
  NAND2X1 U3261 ( .A(arr[1591]), .B(n2671), .Y(n6170) );
  OAI21X1 U3262 ( .A(n4483), .B(n2670), .C(n6171), .Y(n8350) );
  NAND2X1 U3263 ( .A(arr[1592]), .B(n2671), .Y(n6171) );
  OAI21X1 U3264 ( .A(n4485), .B(n2671), .C(n6172), .Y(n8351) );
  NAND2X1 U3265 ( .A(arr[1593]), .B(n2672), .Y(n6172) );
  OAI21X1 U3266 ( .A(n4487), .B(n2671), .C(n6173), .Y(n8352) );
  NAND2X1 U3267 ( .A(arr[1594]), .B(n2672), .Y(n6173) );
  OAI21X1 U3268 ( .A(n4489), .B(n2670), .C(n6174), .Y(n8353) );
  NAND2X1 U3269 ( .A(arr[1595]), .B(n2672), .Y(n6174) );
  OAI21X1 U3270 ( .A(n4491), .B(n2671), .C(n6175), .Y(n8354) );
  NAND2X1 U3271 ( .A(arr[1596]), .B(n2672), .Y(n6175) );
  OAI21X1 U3272 ( .A(n4493), .B(n2671), .C(n6176), .Y(n8355) );
  NAND2X1 U3273 ( .A(arr[1597]), .B(n2672), .Y(n6176) );
  OAI21X1 U3274 ( .A(n4495), .B(n2670), .C(n6177), .Y(n8356) );
  NAND2X1 U3275 ( .A(arr[1598]), .B(n2672), .Y(n6177) );
  OAI21X1 U3276 ( .A(n4497), .B(n2671), .C(n6178), .Y(n8357) );
  NAND2X1 U3277 ( .A(arr[1599]), .B(n2672), .Y(n6178) );
  OAI21X1 U3278 ( .A(n4499), .B(n2671), .C(n6179), .Y(n8358) );
  NAND2X1 U3279 ( .A(arr[1600]), .B(n2672), .Y(n6179) );
  OAI21X1 U3280 ( .A(n4501), .B(n2670), .C(n6180), .Y(n8359) );
  NAND2X1 U3281 ( .A(arr[1601]), .B(n2672), .Y(n6180) );
  OAI21X1 U3282 ( .A(n4503), .B(n2670), .C(n6181), .Y(n8360) );
  NAND2X1 U3283 ( .A(arr[1602]), .B(n2672), .Y(n6181) );
  OAI21X1 U3284 ( .A(n4505), .B(n2670), .C(n6182), .Y(n8361) );
  NAND2X1 U3285 ( .A(arr[1603]), .B(n2672), .Y(n6182) );
  OAI21X1 U3286 ( .A(n4507), .B(n2670), .C(n6183), .Y(n8362) );
  NAND2X1 U3287 ( .A(arr[1604]), .B(n2672), .Y(n6183) );
  OAI21X1 U3288 ( .A(n4509), .B(n2670), .C(n6184), .Y(n8363) );
  NAND2X1 U3289 ( .A(arr[1605]), .B(n2672), .Y(n6184) );
  OAI21X1 U3290 ( .A(n4511), .B(n2670), .C(n6185), .Y(n8364) );
  NAND2X1 U3291 ( .A(arr[1606]), .B(n2672), .Y(n6185) );
  OAI21X1 U3292 ( .A(n4513), .B(n2672), .C(n6186), .Y(n8365) );
  NAND2X1 U3293 ( .A(arr[1607]), .B(n2672), .Y(n6186) );
  OAI21X1 U3294 ( .A(n4515), .B(n2670), .C(n6187), .Y(n8366) );
  NAND2X1 U3295 ( .A(arr[1608]), .B(n2672), .Y(n6187) );
  OAI21X1 U3296 ( .A(n4517), .B(n2671), .C(n6188), .Y(n8367) );
  NAND2X1 U3297 ( .A(arr[1609]), .B(n2672), .Y(n6188) );
  OAI21X1 U3298 ( .A(n4519), .B(n2670), .C(n6189), .Y(n8368) );
  NAND2X1 U3299 ( .A(arr[1610]), .B(n2671), .Y(n6189) );
  OAI21X1 U3300 ( .A(n4521), .B(n2671), .C(n6190), .Y(n8369) );
  NAND2X1 U3301 ( .A(arr[1611]), .B(n2672), .Y(n6190) );
  OAI21X1 U3302 ( .A(n4523), .B(n2670), .C(n6191), .Y(n8370) );
  NAND2X1 U3303 ( .A(arr[1612]), .B(n2671), .Y(n6191) );
  OAI21X1 U3304 ( .A(n4525), .B(n2670), .C(n6192), .Y(n8371) );
  NAND2X1 U3305 ( .A(arr[1613]), .B(n2672), .Y(n6192) );
  OAI21X1 U3306 ( .A(n4527), .B(n2670), .C(n6193), .Y(n8372) );
  NAND2X1 U3307 ( .A(arr[1614]), .B(n2671), .Y(n6193) );
  OAI21X1 U3308 ( .A(n4529), .B(n2670), .C(n6194), .Y(n8373) );
  NAND2X1 U3309 ( .A(arr[1615]), .B(n2671), .Y(n6194) );
  OAI21X1 U3310 ( .A(n4531), .B(n2670), .C(n6195), .Y(n8374) );
  NAND2X1 U3311 ( .A(arr[1616]), .B(n2672), .Y(n6195) );
  OAI21X1 U3313 ( .A(n4467), .B(n2669), .C(n6197), .Y(n8375) );
  NAND2X1 U3314 ( .A(arr[1617]), .B(n2668), .Y(n6197) );
  OAI21X1 U3315 ( .A(n4469), .B(n2667), .C(n6198), .Y(n8376) );
  NAND2X1 U3316 ( .A(arr[1618]), .B(n2668), .Y(n6198) );
  OAI21X1 U3317 ( .A(n4471), .B(n2667), .C(n6199), .Y(n8377) );
  NAND2X1 U3318 ( .A(arr[1619]), .B(n2668), .Y(n6199) );
  OAI21X1 U3319 ( .A(n4473), .B(n2667), .C(n6200), .Y(n8378) );
  NAND2X1 U3320 ( .A(arr[1620]), .B(n2668), .Y(n6200) );
  OAI21X1 U3321 ( .A(n4475), .B(n2667), .C(n6201), .Y(n8379) );
  NAND2X1 U3322 ( .A(arr[1621]), .B(n2668), .Y(n6201) );
  OAI21X1 U3323 ( .A(n4477), .B(n2667), .C(n6202), .Y(n8380) );
  NAND2X1 U3324 ( .A(arr[1622]), .B(n2669), .Y(n6202) );
  OAI21X1 U3325 ( .A(n4479), .B(n2667), .C(n6203), .Y(n8381) );
  NAND2X1 U3326 ( .A(arr[1623]), .B(n2669), .Y(n6203) );
  OAI21X1 U3327 ( .A(n4481), .B(n2668), .C(n6204), .Y(n8382) );
  NAND2X1 U3328 ( .A(arr[1624]), .B(n2668), .Y(n6204) );
  OAI21X1 U3329 ( .A(n4483), .B(n2667), .C(n6205), .Y(n8383) );
  NAND2X1 U3330 ( .A(arr[1625]), .B(n2668), .Y(n6205) );
  OAI21X1 U3331 ( .A(n4485), .B(n2668), .C(n6206), .Y(n8384) );
  NAND2X1 U3332 ( .A(arr[1626]), .B(n2669), .Y(n6206) );
  OAI21X1 U3333 ( .A(n4487), .B(n2668), .C(n6207), .Y(n8385) );
  NAND2X1 U3334 ( .A(arr[1627]), .B(n2669), .Y(n6207) );
  OAI21X1 U3335 ( .A(n4489), .B(n2667), .C(n6208), .Y(n8386) );
  NAND2X1 U3336 ( .A(arr[1628]), .B(n2669), .Y(n6208) );
  OAI21X1 U3337 ( .A(n4491), .B(n2668), .C(n6209), .Y(n8387) );
  NAND2X1 U3338 ( .A(arr[1629]), .B(n2669), .Y(n6209) );
  OAI21X1 U3339 ( .A(n4493), .B(n2668), .C(n6210), .Y(n8388) );
  NAND2X1 U3340 ( .A(arr[1630]), .B(n2669), .Y(n6210) );
  OAI21X1 U3341 ( .A(n4495), .B(n2667), .C(n6211), .Y(n8389) );
  NAND2X1 U3342 ( .A(arr[1631]), .B(n2669), .Y(n6211) );
  OAI21X1 U3343 ( .A(n4497), .B(n2668), .C(n6212), .Y(n8390) );
  NAND2X1 U3344 ( .A(arr[1632]), .B(n2669), .Y(n6212) );
  OAI21X1 U3345 ( .A(n4499), .B(n2668), .C(n6213), .Y(n8391) );
  NAND2X1 U3346 ( .A(arr[1633]), .B(n2669), .Y(n6213) );
  OAI21X1 U3347 ( .A(n4501), .B(n2667), .C(n6214), .Y(n8392) );
  NAND2X1 U3348 ( .A(arr[1634]), .B(n2669), .Y(n6214) );
  OAI21X1 U3349 ( .A(n4503), .B(n2667), .C(n6215), .Y(n8393) );
  NAND2X1 U3350 ( .A(arr[1635]), .B(n2669), .Y(n6215) );
  OAI21X1 U3351 ( .A(n4505), .B(n2667), .C(n6216), .Y(n8394) );
  NAND2X1 U3352 ( .A(arr[1636]), .B(n2669), .Y(n6216) );
  OAI21X1 U3353 ( .A(n4507), .B(n2667), .C(n6217), .Y(n8395) );
  NAND2X1 U3354 ( .A(arr[1637]), .B(n2669), .Y(n6217) );
  OAI21X1 U3355 ( .A(n4509), .B(n2667), .C(n6218), .Y(n8396) );
  NAND2X1 U3356 ( .A(arr[1638]), .B(n2669), .Y(n6218) );
  OAI21X1 U3357 ( .A(n4511), .B(n2667), .C(n6219), .Y(n8397) );
  NAND2X1 U3358 ( .A(arr[1639]), .B(n2669), .Y(n6219) );
  OAI21X1 U3359 ( .A(n4513), .B(n2669), .C(n6220), .Y(n8398) );
  NAND2X1 U3360 ( .A(arr[1640]), .B(n2669), .Y(n6220) );
  OAI21X1 U3361 ( .A(n4515), .B(n2667), .C(n6221), .Y(n8399) );
  NAND2X1 U3362 ( .A(arr[1641]), .B(n2669), .Y(n6221) );
  OAI21X1 U3363 ( .A(n4517), .B(n2668), .C(n6222), .Y(n8400) );
  NAND2X1 U3364 ( .A(arr[1642]), .B(n2669), .Y(n6222) );
  OAI21X1 U3365 ( .A(n4519), .B(n2667), .C(n6223), .Y(n8401) );
  NAND2X1 U3366 ( .A(arr[1643]), .B(n2668), .Y(n6223) );
  OAI21X1 U3367 ( .A(n4521), .B(n2668), .C(n6224), .Y(n8402) );
  NAND2X1 U3368 ( .A(arr[1644]), .B(n2669), .Y(n6224) );
  OAI21X1 U3369 ( .A(n4523), .B(n2667), .C(n6225), .Y(n8403) );
  NAND2X1 U3370 ( .A(arr[1645]), .B(n2668), .Y(n6225) );
  OAI21X1 U3371 ( .A(n4525), .B(n2667), .C(n6226), .Y(n8404) );
  NAND2X1 U3372 ( .A(arr[1646]), .B(n2669), .Y(n6226) );
  OAI21X1 U3373 ( .A(n4527), .B(n2667), .C(n6227), .Y(n8405) );
  NAND2X1 U3374 ( .A(arr[1647]), .B(n2668), .Y(n6227) );
  OAI21X1 U3375 ( .A(n4529), .B(n2667), .C(n6228), .Y(n8406) );
  NAND2X1 U3376 ( .A(arr[1648]), .B(n2668), .Y(n6228) );
  OAI21X1 U3377 ( .A(n4531), .B(n2667), .C(n6229), .Y(n8407) );
  NAND2X1 U3378 ( .A(arr[1649]), .B(n2669), .Y(n6229) );
  AND2X1 U3380 ( .A(n6230), .B(n5680), .Y(n5087) );
  OAI21X1 U3381 ( .A(n4467), .B(n2666), .C(n6232), .Y(n8408) );
  NAND2X1 U3382 ( .A(arr[1650]), .B(n2665), .Y(n6232) );
  OAI21X1 U3383 ( .A(n4469), .B(n2664), .C(n6233), .Y(n8409) );
  NAND2X1 U3384 ( .A(arr[1651]), .B(n2665), .Y(n6233) );
  OAI21X1 U3385 ( .A(n4471), .B(n2664), .C(n6234), .Y(n8410) );
  NAND2X1 U3386 ( .A(arr[1652]), .B(n2665), .Y(n6234) );
  OAI21X1 U3387 ( .A(n4473), .B(n2664), .C(n6235), .Y(n8411) );
  NAND2X1 U3388 ( .A(arr[1653]), .B(n2665), .Y(n6235) );
  OAI21X1 U3389 ( .A(n4475), .B(n2664), .C(n6236), .Y(n8412) );
  NAND2X1 U3390 ( .A(arr[1654]), .B(n2665), .Y(n6236) );
  OAI21X1 U3391 ( .A(n4477), .B(n2664), .C(n6237), .Y(n8413) );
  NAND2X1 U3392 ( .A(arr[1655]), .B(n2666), .Y(n6237) );
  OAI21X1 U3393 ( .A(n4479), .B(n2664), .C(n6238), .Y(n8414) );
  NAND2X1 U3394 ( .A(arr[1656]), .B(n2666), .Y(n6238) );
  OAI21X1 U3395 ( .A(n4481), .B(n2665), .C(n6239), .Y(n8415) );
  NAND2X1 U3396 ( .A(arr[1657]), .B(n2665), .Y(n6239) );
  OAI21X1 U3397 ( .A(n4483), .B(n2664), .C(n6240), .Y(n8416) );
  NAND2X1 U3398 ( .A(arr[1658]), .B(n2665), .Y(n6240) );
  OAI21X1 U3399 ( .A(n4485), .B(n2665), .C(n6241), .Y(n8417) );
  NAND2X1 U3400 ( .A(arr[1659]), .B(n2666), .Y(n6241) );
  OAI21X1 U3401 ( .A(n4487), .B(n2665), .C(n6242), .Y(n8418) );
  NAND2X1 U3402 ( .A(arr[1660]), .B(n2666), .Y(n6242) );
  OAI21X1 U3403 ( .A(n4489), .B(n2664), .C(n6243), .Y(n8419) );
  NAND2X1 U3404 ( .A(arr[1661]), .B(n2666), .Y(n6243) );
  OAI21X1 U3405 ( .A(n4491), .B(n2665), .C(n6244), .Y(n8420) );
  NAND2X1 U3406 ( .A(arr[1662]), .B(n2666), .Y(n6244) );
  OAI21X1 U3407 ( .A(n4493), .B(n2665), .C(n6245), .Y(n8421) );
  NAND2X1 U3408 ( .A(arr[1663]), .B(n2666), .Y(n6245) );
  OAI21X1 U3409 ( .A(n4495), .B(n2664), .C(n6246), .Y(n8422) );
  NAND2X1 U3410 ( .A(arr[1664]), .B(n2666), .Y(n6246) );
  OAI21X1 U3411 ( .A(n4497), .B(n2665), .C(n6247), .Y(n8423) );
  NAND2X1 U3412 ( .A(arr[1665]), .B(n2666), .Y(n6247) );
  OAI21X1 U3413 ( .A(n4499), .B(n2665), .C(n6248), .Y(n8424) );
  NAND2X1 U3414 ( .A(arr[1666]), .B(n2666), .Y(n6248) );
  OAI21X1 U3415 ( .A(n4501), .B(n2664), .C(n6249), .Y(n8425) );
  NAND2X1 U3416 ( .A(arr[1667]), .B(n2666), .Y(n6249) );
  OAI21X1 U3417 ( .A(n4503), .B(n2664), .C(n6250), .Y(n8426) );
  NAND2X1 U3418 ( .A(arr[1668]), .B(n2666), .Y(n6250) );
  OAI21X1 U3419 ( .A(n4505), .B(n2664), .C(n6251), .Y(n8427) );
  NAND2X1 U3420 ( .A(arr[1669]), .B(n2666), .Y(n6251) );
  OAI21X1 U3421 ( .A(n4507), .B(n2664), .C(n6252), .Y(n8428) );
  NAND2X1 U3422 ( .A(arr[1670]), .B(n2666), .Y(n6252) );
  OAI21X1 U3423 ( .A(n4509), .B(n2664), .C(n6253), .Y(n8429) );
  NAND2X1 U3424 ( .A(arr[1671]), .B(n2666), .Y(n6253) );
  OAI21X1 U3425 ( .A(n4511), .B(n2664), .C(n6254), .Y(n8430) );
  NAND2X1 U3426 ( .A(arr[1672]), .B(n2666), .Y(n6254) );
  OAI21X1 U3427 ( .A(n4513), .B(n2666), .C(n6255), .Y(n8431) );
  NAND2X1 U3428 ( .A(arr[1673]), .B(n2666), .Y(n6255) );
  OAI21X1 U3429 ( .A(n4515), .B(n2664), .C(n6256), .Y(n8432) );
  NAND2X1 U3430 ( .A(arr[1674]), .B(n2666), .Y(n6256) );
  OAI21X1 U3431 ( .A(n4517), .B(n2665), .C(n6257), .Y(n8433) );
  NAND2X1 U3432 ( .A(arr[1675]), .B(n2666), .Y(n6257) );
  OAI21X1 U3433 ( .A(n4519), .B(n2664), .C(n6258), .Y(n8434) );
  NAND2X1 U3434 ( .A(arr[1676]), .B(n2665), .Y(n6258) );
  OAI21X1 U3435 ( .A(n4521), .B(n2665), .C(n6259), .Y(n8435) );
  NAND2X1 U3436 ( .A(arr[1677]), .B(n2666), .Y(n6259) );
  OAI21X1 U3437 ( .A(n4523), .B(n2664), .C(n6260), .Y(n8436) );
  NAND2X1 U3438 ( .A(arr[1678]), .B(n2665), .Y(n6260) );
  OAI21X1 U3439 ( .A(n4525), .B(n2664), .C(n6261), .Y(n8437) );
  NAND2X1 U3440 ( .A(arr[1679]), .B(n2666), .Y(n6261) );
  OAI21X1 U3441 ( .A(n4527), .B(n2664), .C(n6262), .Y(n8438) );
  NAND2X1 U3442 ( .A(arr[1680]), .B(n2665), .Y(n6262) );
  OAI21X1 U3443 ( .A(n4529), .B(n2664), .C(n6263), .Y(n8439) );
  NAND2X1 U3444 ( .A(arr[1681]), .B(n2665), .Y(n6263) );
  OAI21X1 U3445 ( .A(n4531), .B(n2664), .C(n6264), .Y(n8440) );
  NAND2X1 U3446 ( .A(arr[1682]), .B(n2666), .Y(n6264) );
  OAI21X1 U3448 ( .A(n4467), .B(n2663), .C(n6266), .Y(n8441) );
  NAND2X1 U3449 ( .A(arr[1683]), .B(n2662), .Y(n6266) );
  OAI21X1 U3450 ( .A(n4469), .B(n2661), .C(n6267), .Y(n8442) );
  NAND2X1 U3451 ( .A(arr[1684]), .B(n2662), .Y(n6267) );
  OAI21X1 U3452 ( .A(n4471), .B(n2661), .C(n6268), .Y(n8443) );
  NAND2X1 U3453 ( .A(arr[1685]), .B(n2662), .Y(n6268) );
  OAI21X1 U3454 ( .A(n4473), .B(n2661), .C(n6269), .Y(n8444) );
  NAND2X1 U3455 ( .A(arr[1686]), .B(n2662), .Y(n6269) );
  OAI21X1 U3456 ( .A(n4475), .B(n2661), .C(n6270), .Y(n8445) );
  NAND2X1 U3457 ( .A(arr[1687]), .B(n2662), .Y(n6270) );
  OAI21X1 U3458 ( .A(n4477), .B(n2661), .C(n6271), .Y(n8446) );
  NAND2X1 U3459 ( .A(arr[1688]), .B(n2663), .Y(n6271) );
  OAI21X1 U3460 ( .A(n4479), .B(n2661), .C(n6272), .Y(n8447) );
  NAND2X1 U3461 ( .A(arr[1689]), .B(n2663), .Y(n6272) );
  OAI21X1 U3462 ( .A(n4481), .B(n2662), .C(n6273), .Y(n8448) );
  NAND2X1 U3463 ( .A(arr[1690]), .B(n2662), .Y(n6273) );
  OAI21X1 U3464 ( .A(n4483), .B(n2661), .C(n6274), .Y(n8449) );
  NAND2X1 U3465 ( .A(arr[1691]), .B(n2662), .Y(n6274) );
  OAI21X1 U3466 ( .A(n4485), .B(n2662), .C(n6275), .Y(n8450) );
  NAND2X1 U3467 ( .A(arr[1692]), .B(n2663), .Y(n6275) );
  OAI21X1 U3468 ( .A(n4487), .B(n2662), .C(n6276), .Y(n8451) );
  NAND2X1 U3469 ( .A(arr[1693]), .B(n2663), .Y(n6276) );
  OAI21X1 U3470 ( .A(n4489), .B(n2661), .C(n6277), .Y(n8452) );
  NAND2X1 U3471 ( .A(arr[1694]), .B(n2663), .Y(n6277) );
  OAI21X1 U3472 ( .A(n4491), .B(n2662), .C(n6278), .Y(n8453) );
  NAND2X1 U3473 ( .A(arr[1695]), .B(n2663), .Y(n6278) );
  OAI21X1 U3474 ( .A(n4493), .B(n2662), .C(n6279), .Y(n8454) );
  NAND2X1 U3475 ( .A(arr[1696]), .B(n2663), .Y(n6279) );
  OAI21X1 U3476 ( .A(n4495), .B(n2661), .C(n6280), .Y(n8455) );
  NAND2X1 U3477 ( .A(arr[1697]), .B(n2663), .Y(n6280) );
  OAI21X1 U3478 ( .A(n4497), .B(n2662), .C(n6281), .Y(n8456) );
  NAND2X1 U3479 ( .A(arr[1698]), .B(n2663), .Y(n6281) );
  OAI21X1 U3480 ( .A(n4499), .B(n2662), .C(n6282), .Y(n8457) );
  NAND2X1 U3481 ( .A(arr[1699]), .B(n2663), .Y(n6282) );
  OAI21X1 U3482 ( .A(n4501), .B(n2661), .C(n6283), .Y(n8458) );
  NAND2X1 U3483 ( .A(arr[1700]), .B(n2663), .Y(n6283) );
  OAI21X1 U3484 ( .A(n4503), .B(n2661), .C(n6284), .Y(n8459) );
  NAND2X1 U3485 ( .A(arr[1701]), .B(n2663), .Y(n6284) );
  OAI21X1 U3486 ( .A(n4505), .B(n2661), .C(n6285), .Y(n8460) );
  NAND2X1 U3487 ( .A(arr[1702]), .B(n2663), .Y(n6285) );
  OAI21X1 U3488 ( .A(n4507), .B(n2661), .C(n6286), .Y(n8461) );
  NAND2X1 U3489 ( .A(arr[1703]), .B(n2663), .Y(n6286) );
  OAI21X1 U3490 ( .A(n4509), .B(n2661), .C(n6287), .Y(n8462) );
  NAND2X1 U3491 ( .A(arr[1704]), .B(n2663), .Y(n6287) );
  OAI21X1 U3492 ( .A(n4511), .B(n2661), .C(n6288), .Y(n8463) );
  NAND2X1 U3493 ( .A(arr[1705]), .B(n2663), .Y(n6288) );
  OAI21X1 U3494 ( .A(n4513), .B(n2663), .C(n6289), .Y(n8464) );
  NAND2X1 U3495 ( .A(arr[1706]), .B(n2663), .Y(n6289) );
  OAI21X1 U3496 ( .A(n4515), .B(n2661), .C(n6290), .Y(n8465) );
  NAND2X1 U3497 ( .A(arr[1707]), .B(n2663), .Y(n6290) );
  OAI21X1 U3498 ( .A(n4517), .B(n2662), .C(n6291), .Y(n8466) );
  NAND2X1 U3499 ( .A(arr[1708]), .B(n2663), .Y(n6291) );
  OAI21X1 U3500 ( .A(n4519), .B(n2661), .C(n6292), .Y(n8467) );
  NAND2X1 U3501 ( .A(arr[1709]), .B(n2662), .Y(n6292) );
  OAI21X1 U3502 ( .A(n4521), .B(n2662), .C(n6293), .Y(n8468) );
  NAND2X1 U3503 ( .A(arr[1710]), .B(n2663), .Y(n6293) );
  OAI21X1 U3504 ( .A(n4523), .B(n2661), .C(n6294), .Y(n8469) );
  NAND2X1 U3505 ( .A(arr[1711]), .B(n2662), .Y(n6294) );
  OAI21X1 U3506 ( .A(n4525), .B(n2661), .C(n6295), .Y(n8470) );
  NAND2X1 U3507 ( .A(arr[1712]), .B(n2663), .Y(n6295) );
  OAI21X1 U3508 ( .A(n4527), .B(n2661), .C(n6296), .Y(n8471) );
  NAND2X1 U3509 ( .A(arr[1713]), .B(n2662), .Y(n6296) );
  OAI21X1 U3510 ( .A(n4529), .B(n2661), .C(n6297), .Y(n8472) );
  NAND2X1 U3511 ( .A(arr[1714]), .B(n2662), .Y(n6297) );
  OAI21X1 U3512 ( .A(n4531), .B(n2661), .C(n6298), .Y(n8473) );
  NAND2X1 U3513 ( .A(arr[1715]), .B(n2663), .Y(n6298) );
  AND2X1 U3515 ( .A(n6230), .B(n5749), .Y(n5156) );
  OAI21X1 U3516 ( .A(n4467), .B(n2660), .C(n6300), .Y(n8474) );
  NAND2X1 U3517 ( .A(arr[1716]), .B(n2659), .Y(n6300) );
  OAI21X1 U3518 ( .A(n4469), .B(n2658), .C(n6301), .Y(n8475) );
  NAND2X1 U3519 ( .A(arr[1717]), .B(n2659), .Y(n6301) );
  OAI21X1 U3520 ( .A(n4471), .B(n2658), .C(n6302), .Y(n8476) );
  NAND2X1 U3521 ( .A(arr[1718]), .B(n2659), .Y(n6302) );
  OAI21X1 U3522 ( .A(n4473), .B(n2658), .C(n6303), .Y(n8477) );
  NAND2X1 U3523 ( .A(arr[1719]), .B(n2659), .Y(n6303) );
  OAI21X1 U3524 ( .A(n4475), .B(n2658), .C(n6304), .Y(n8478) );
  NAND2X1 U3525 ( .A(arr[1720]), .B(n2659), .Y(n6304) );
  OAI21X1 U3526 ( .A(n4477), .B(n2658), .C(n6305), .Y(n8479) );
  NAND2X1 U3527 ( .A(arr[1721]), .B(n2660), .Y(n6305) );
  OAI21X1 U3528 ( .A(n4479), .B(n2658), .C(n6306), .Y(n8480) );
  NAND2X1 U3529 ( .A(arr[1722]), .B(n2660), .Y(n6306) );
  OAI21X1 U3530 ( .A(n4481), .B(n2659), .C(n6307), .Y(n8481) );
  NAND2X1 U3531 ( .A(arr[1723]), .B(n2659), .Y(n6307) );
  OAI21X1 U3532 ( .A(n4483), .B(n2658), .C(n6308), .Y(n8482) );
  NAND2X1 U3533 ( .A(arr[1724]), .B(n2659), .Y(n6308) );
  OAI21X1 U3534 ( .A(n4485), .B(n2659), .C(n6309), .Y(n8483) );
  NAND2X1 U3535 ( .A(arr[1725]), .B(n2660), .Y(n6309) );
  OAI21X1 U3536 ( .A(n4487), .B(n2659), .C(n6310), .Y(n8484) );
  NAND2X1 U3537 ( .A(arr[1726]), .B(n2660), .Y(n6310) );
  OAI21X1 U3538 ( .A(n4489), .B(n2658), .C(n6311), .Y(n8485) );
  NAND2X1 U3539 ( .A(arr[1727]), .B(n2660), .Y(n6311) );
  OAI21X1 U3540 ( .A(n4491), .B(n2659), .C(n6312), .Y(n8486) );
  NAND2X1 U3541 ( .A(arr[1728]), .B(n2660), .Y(n6312) );
  OAI21X1 U3542 ( .A(n4493), .B(n2659), .C(n6313), .Y(n8487) );
  NAND2X1 U3543 ( .A(arr[1729]), .B(n2660), .Y(n6313) );
  OAI21X1 U3544 ( .A(n4495), .B(n2658), .C(n6314), .Y(n8488) );
  NAND2X1 U3545 ( .A(arr[1730]), .B(n2660), .Y(n6314) );
  OAI21X1 U3546 ( .A(n4497), .B(n2659), .C(n6315), .Y(n8489) );
  NAND2X1 U3547 ( .A(arr[1731]), .B(n2660), .Y(n6315) );
  OAI21X1 U3548 ( .A(n4499), .B(n2659), .C(n6316), .Y(n8490) );
  NAND2X1 U3549 ( .A(arr[1732]), .B(n2660), .Y(n6316) );
  OAI21X1 U3550 ( .A(n4501), .B(n2658), .C(n6317), .Y(n8491) );
  NAND2X1 U3551 ( .A(arr[1733]), .B(n2660), .Y(n6317) );
  OAI21X1 U3552 ( .A(n4503), .B(n2658), .C(n6318), .Y(n8492) );
  NAND2X1 U3553 ( .A(arr[1734]), .B(n2660), .Y(n6318) );
  OAI21X1 U3554 ( .A(n4505), .B(n2658), .C(n6319), .Y(n8493) );
  NAND2X1 U3555 ( .A(arr[1735]), .B(n2660), .Y(n6319) );
  OAI21X1 U3556 ( .A(n4507), .B(n2658), .C(n6320), .Y(n8494) );
  NAND2X1 U3557 ( .A(arr[1736]), .B(n2660), .Y(n6320) );
  OAI21X1 U3558 ( .A(n4509), .B(n2658), .C(n6321), .Y(n8495) );
  NAND2X1 U3559 ( .A(arr[1737]), .B(n2660), .Y(n6321) );
  OAI21X1 U3560 ( .A(n4511), .B(n2658), .C(n6322), .Y(n8496) );
  NAND2X1 U3561 ( .A(arr[1738]), .B(n2660), .Y(n6322) );
  OAI21X1 U3562 ( .A(n4513), .B(n2660), .C(n6323), .Y(n8497) );
  NAND2X1 U3563 ( .A(arr[1739]), .B(n2660), .Y(n6323) );
  OAI21X1 U3564 ( .A(n4515), .B(n2658), .C(n6324), .Y(n8498) );
  NAND2X1 U3565 ( .A(arr[1740]), .B(n2660), .Y(n6324) );
  OAI21X1 U3566 ( .A(n4517), .B(n2659), .C(n6325), .Y(n8499) );
  NAND2X1 U3567 ( .A(arr[1741]), .B(n2660), .Y(n6325) );
  OAI21X1 U3568 ( .A(n4519), .B(n2658), .C(n6326), .Y(n8500) );
  NAND2X1 U3569 ( .A(arr[1742]), .B(n2659), .Y(n6326) );
  OAI21X1 U3570 ( .A(n4521), .B(n2659), .C(n6327), .Y(n8501) );
  NAND2X1 U3571 ( .A(arr[1743]), .B(n2660), .Y(n6327) );
  OAI21X1 U3572 ( .A(n4523), .B(n2658), .C(n6328), .Y(n8502) );
  NAND2X1 U3573 ( .A(arr[1744]), .B(n2659), .Y(n6328) );
  OAI21X1 U3574 ( .A(n4525), .B(n2658), .C(n6329), .Y(n8503) );
  NAND2X1 U3575 ( .A(arr[1745]), .B(n2660), .Y(n6329) );
  OAI21X1 U3576 ( .A(n4527), .B(n2658), .C(n6330), .Y(n8504) );
  NAND2X1 U3577 ( .A(arr[1746]), .B(n2659), .Y(n6330) );
  OAI21X1 U3578 ( .A(n4529), .B(n2658), .C(n6331), .Y(n8505) );
  NAND2X1 U3579 ( .A(arr[1747]), .B(n2659), .Y(n6331) );
  OAI21X1 U3580 ( .A(n4531), .B(n2658), .C(n6332), .Y(n8506) );
  NAND2X1 U3581 ( .A(arr[1748]), .B(n2660), .Y(n6332) );
  OAI21X1 U3583 ( .A(n4467), .B(n2657), .C(n6334), .Y(n8507) );
  NAND2X1 U3584 ( .A(arr[1749]), .B(n2656), .Y(n6334) );
  OAI21X1 U3585 ( .A(n4469), .B(n2655), .C(n6335), .Y(n8508) );
  NAND2X1 U3586 ( .A(arr[1750]), .B(n2656), .Y(n6335) );
  OAI21X1 U3587 ( .A(n4471), .B(n2655), .C(n6336), .Y(n8509) );
  NAND2X1 U3588 ( .A(arr[1751]), .B(n2656), .Y(n6336) );
  OAI21X1 U3589 ( .A(n4473), .B(n2655), .C(n6337), .Y(n8510) );
  NAND2X1 U3590 ( .A(arr[1752]), .B(n2656), .Y(n6337) );
  OAI21X1 U3591 ( .A(n4475), .B(n2655), .C(n6338), .Y(n8511) );
  NAND2X1 U3592 ( .A(arr[1753]), .B(n2656), .Y(n6338) );
  OAI21X1 U3593 ( .A(n4477), .B(n2655), .C(n6339), .Y(n8512) );
  NAND2X1 U3594 ( .A(arr[1754]), .B(n2657), .Y(n6339) );
  OAI21X1 U3595 ( .A(n4479), .B(n2655), .C(n6340), .Y(n8513) );
  NAND2X1 U3596 ( .A(arr[1755]), .B(n2657), .Y(n6340) );
  OAI21X1 U3597 ( .A(n4481), .B(n2656), .C(n6341), .Y(n8514) );
  NAND2X1 U3598 ( .A(arr[1756]), .B(n2656), .Y(n6341) );
  OAI21X1 U3599 ( .A(n4483), .B(n2655), .C(n6342), .Y(n8515) );
  NAND2X1 U3600 ( .A(arr[1757]), .B(n2656), .Y(n6342) );
  OAI21X1 U3601 ( .A(n4485), .B(n2656), .C(n6343), .Y(n8516) );
  NAND2X1 U3602 ( .A(arr[1758]), .B(n2657), .Y(n6343) );
  OAI21X1 U3603 ( .A(n4487), .B(n2656), .C(n6344), .Y(n8517) );
  NAND2X1 U3604 ( .A(arr[1759]), .B(n2657), .Y(n6344) );
  OAI21X1 U3605 ( .A(n4489), .B(n2655), .C(n6345), .Y(n8518) );
  NAND2X1 U3606 ( .A(arr[1760]), .B(n2657), .Y(n6345) );
  OAI21X1 U3607 ( .A(n4491), .B(n2656), .C(n6346), .Y(n8519) );
  NAND2X1 U3608 ( .A(arr[1761]), .B(n2657), .Y(n6346) );
  OAI21X1 U3609 ( .A(n4493), .B(n2656), .C(n6347), .Y(n8520) );
  NAND2X1 U3610 ( .A(arr[1762]), .B(n2657), .Y(n6347) );
  OAI21X1 U3611 ( .A(n4495), .B(n2655), .C(n6348), .Y(n8521) );
  NAND2X1 U3612 ( .A(arr[1763]), .B(n2657), .Y(n6348) );
  OAI21X1 U3613 ( .A(n4497), .B(n2656), .C(n6349), .Y(n8522) );
  NAND2X1 U3614 ( .A(arr[1764]), .B(n2657), .Y(n6349) );
  OAI21X1 U3615 ( .A(n4499), .B(n2656), .C(n6350), .Y(n8523) );
  NAND2X1 U3616 ( .A(arr[1765]), .B(n2657), .Y(n6350) );
  OAI21X1 U3617 ( .A(n4501), .B(n2655), .C(n6351), .Y(n8524) );
  NAND2X1 U3618 ( .A(arr[1766]), .B(n2657), .Y(n6351) );
  OAI21X1 U3619 ( .A(n4503), .B(n2655), .C(n6352), .Y(n8525) );
  NAND2X1 U3620 ( .A(arr[1767]), .B(n2657), .Y(n6352) );
  OAI21X1 U3621 ( .A(n4505), .B(n2655), .C(n6353), .Y(n8526) );
  NAND2X1 U3622 ( .A(arr[1768]), .B(n2657), .Y(n6353) );
  OAI21X1 U3623 ( .A(n4507), .B(n2655), .C(n6354), .Y(n8527) );
  NAND2X1 U3624 ( .A(arr[1769]), .B(n2657), .Y(n6354) );
  OAI21X1 U3625 ( .A(n4509), .B(n2655), .C(n6355), .Y(n8528) );
  NAND2X1 U3626 ( .A(arr[1770]), .B(n2657), .Y(n6355) );
  OAI21X1 U3627 ( .A(n4511), .B(n2655), .C(n6356), .Y(n8529) );
  NAND2X1 U3628 ( .A(arr[1771]), .B(n2657), .Y(n6356) );
  OAI21X1 U3629 ( .A(n4513), .B(n2657), .C(n6357), .Y(n8530) );
  NAND2X1 U3630 ( .A(arr[1772]), .B(n2657), .Y(n6357) );
  OAI21X1 U3631 ( .A(n4515), .B(n2655), .C(n6358), .Y(n8531) );
  NAND2X1 U3632 ( .A(arr[1773]), .B(n2657), .Y(n6358) );
  OAI21X1 U3633 ( .A(n4517), .B(n2656), .C(n6359), .Y(n8532) );
  NAND2X1 U3634 ( .A(arr[1774]), .B(n2657), .Y(n6359) );
  OAI21X1 U3635 ( .A(n4519), .B(n2655), .C(n6360), .Y(n8533) );
  NAND2X1 U3636 ( .A(arr[1775]), .B(n2656), .Y(n6360) );
  OAI21X1 U3637 ( .A(n4521), .B(n2656), .C(n6361), .Y(n8534) );
  NAND2X1 U3638 ( .A(arr[1776]), .B(n2657), .Y(n6361) );
  OAI21X1 U3639 ( .A(n4523), .B(n2655), .C(n6362), .Y(n8535) );
  NAND2X1 U3640 ( .A(arr[1777]), .B(n2656), .Y(n6362) );
  OAI21X1 U3641 ( .A(n4525), .B(n2655), .C(n6363), .Y(n8536) );
  NAND2X1 U3642 ( .A(arr[1778]), .B(n2657), .Y(n6363) );
  OAI21X1 U3643 ( .A(n4527), .B(n2655), .C(n6364), .Y(n8537) );
  NAND2X1 U3644 ( .A(arr[1779]), .B(n2656), .Y(n6364) );
  OAI21X1 U3645 ( .A(n4529), .B(n2655), .C(n6365), .Y(n8538) );
  NAND2X1 U3646 ( .A(arr[1780]), .B(n2656), .Y(n6365) );
  OAI21X1 U3647 ( .A(n4531), .B(n2655), .C(n6366), .Y(n8539) );
  NAND2X1 U3648 ( .A(arr[1781]), .B(n2657), .Y(n6366) );
  AND2X1 U3650 ( .A(n6230), .B(n5818), .Y(n5225) );
  OAI21X1 U3651 ( .A(n4467), .B(n2654), .C(n6368), .Y(n8540) );
  NAND2X1 U3652 ( .A(arr[1782]), .B(n2653), .Y(n6368) );
  OAI21X1 U3653 ( .A(n4469), .B(n2652), .C(n6369), .Y(n8541) );
  NAND2X1 U3654 ( .A(arr[1783]), .B(n2653), .Y(n6369) );
  OAI21X1 U3655 ( .A(n4471), .B(n2652), .C(n6370), .Y(n8542) );
  NAND2X1 U3656 ( .A(arr[1784]), .B(n2653), .Y(n6370) );
  OAI21X1 U3657 ( .A(n4473), .B(n2652), .C(n6371), .Y(n8543) );
  NAND2X1 U3658 ( .A(arr[1785]), .B(n2653), .Y(n6371) );
  OAI21X1 U3659 ( .A(n4475), .B(n2652), .C(n6372), .Y(n8544) );
  NAND2X1 U3660 ( .A(arr[1786]), .B(n2653), .Y(n6372) );
  OAI21X1 U3661 ( .A(n4477), .B(n2652), .C(n6373), .Y(n8545) );
  NAND2X1 U3662 ( .A(arr[1787]), .B(n2654), .Y(n6373) );
  OAI21X1 U3663 ( .A(n4479), .B(n2652), .C(n6374), .Y(n8546) );
  NAND2X1 U3664 ( .A(arr[1788]), .B(n2654), .Y(n6374) );
  OAI21X1 U3665 ( .A(n4481), .B(n2653), .C(n6375), .Y(n8547) );
  NAND2X1 U3666 ( .A(arr[1789]), .B(n2653), .Y(n6375) );
  OAI21X1 U3667 ( .A(n4483), .B(n2652), .C(n6376), .Y(n8548) );
  NAND2X1 U3668 ( .A(arr[1790]), .B(n2653), .Y(n6376) );
  OAI21X1 U3669 ( .A(n4485), .B(n2653), .C(n6377), .Y(n8549) );
  NAND2X1 U3670 ( .A(arr[1791]), .B(n2654), .Y(n6377) );
  OAI21X1 U3671 ( .A(n4487), .B(n2653), .C(n6378), .Y(n8550) );
  NAND2X1 U3672 ( .A(arr[1792]), .B(n2654), .Y(n6378) );
  OAI21X1 U3673 ( .A(n4489), .B(n2652), .C(n6379), .Y(n8551) );
  NAND2X1 U3674 ( .A(arr[1793]), .B(n2654), .Y(n6379) );
  OAI21X1 U3675 ( .A(n4491), .B(n2653), .C(n6380), .Y(n8552) );
  NAND2X1 U3676 ( .A(arr[1794]), .B(n2654), .Y(n6380) );
  OAI21X1 U3677 ( .A(n4493), .B(n2653), .C(n6381), .Y(n8553) );
  NAND2X1 U3678 ( .A(arr[1795]), .B(n2654), .Y(n6381) );
  OAI21X1 U3679 ( .A(n4495), .B(n2652), .C(n6382), .Y(n8554) );
  NAND2X1 U3680 ( .A(arr[1796]), .B(n2654), .Y(n6382) );
  OAI21X1 U3681 ( .A(n4497), .B(n2653), .C(n6383), .Y(n8555) );
  NAND2X1 U3682 ( .A(arr[1797]), .B(n2654), .Y(n6383) );
  OAI21X1 U3683 ( .A(n4499), .B(n2653), .C(n6384), .Y(n8556) );
  NAND2X1 U3684 ( .A(arr[1798]), .B(n2654), .Y(n6384) );
  OAI21X1 U3685 ( .A(n4501), .B(n2652), .C(n6385), .Y(n8557) );
  NAND2X1 U3686 ( .A(arr[1799]), .B(n2654), .Y(n6385) );
  OAI21X1 U3687 ( .A(n4503), .B(n2652), .C(n6386), .Y(n8558) );
  NAND2X1 U3688 ( .A(arr[1800]), .B(n2654), .Y(n6386) );
  OAI21X1 U3689 ( .A(n4505), .B(n2652), .C(n6387), .Y(n8559) );
  NAND2X1 U3690 ( .A(arr[1801]), .B(n2654), .Y(n6387) );
  OAI21X1 U3691 ( .A(n4507), .B(n2652), .C(n6388), .Y(n8560) );
  NAND2X1 U3692 ( .A(arr[1802]), .B(n2654), .Y(n6388) );
  OAI21X1 U3693 ( .A(n4509), .B(n2652), .C(n6389), .Y(n8561) );
  NAND2X1 U3694 ( .A(arr[1803]), .B(n2654), .Y(n6389) );
  OAI21X1 U3695 ( .A(n4511), .B(n2652), .C(n6390), .Y(n8562) );
  NAND2X1 U3696 ( .A(arr[1804]), .B(n2654), .Y(n6390) );
  OAI21X1 U3697 ( .A(n4513), .B(n2654), .C(n6391), .Y(n8563) );
  NAND2X1 U3698 ( .A(arr[1805]), .B(n2654), .Y(n6391) );
  OAI21X1 U3699 ( .A(n4515), .B(n2652), .C(n6392), .Y(n8564) );
  NAND2X1 U3700 ( .A(arr[1806]), .B(n2654), .Y(n6392) );
  OAI21X1 U3701 ( .A(n4517), .B(n2653), .C(n6393), .Y(n8565) );
  NAND2X1 U3702 ( .A(arr[1807]), .B(n2654), .Y(n6393) );
  OAI21X1 U3703 ( .A(n4519), .B(n2652), .C(n6394), .Y(n8566) );
  NAND2X1 U3704 ( .A(arr[1808]), .B(n2653), .Y(n6394) );
  OAI21X1 U3705 ( .A(n4521), .B(n2653), .C(n6395), .Y(n8567) );
  NAND2X1 U3706 ( .A(arr[1809]), .B(n2654), .Y(n6395) );
  OAI21X1 U3707 ( .A(n4523), .B(n2652), .C(n6396), .Y(n8568) );
  NAND2X1 U3708 ( .A(arr[1810]), .B(n2653), .Y(n6396) );
  OAI21X1 U3709 ( .A(n4525), .B(n2652), .C(n6397), .Y(n8569) );
  NAND2X1 U3710 ( .A(arr[1811]), .B(n2654), .Y(n6397) );
  OAI21X1 U3711 ( .A(n4527), .B(n2652), .C(n6398), .Y(n8570) );
  NAND2X1 U3712 ( .A(arr[1812]), .B(n2653), .Y(n6398) );
  OAI21X1 U3713 ( .A(n4529), .B(n2652), .C(n6399), .Y(n8571) );
  NAND2X1 U3714 ( .A(arr[1813]), .B(n2653), .Y(n6399) );
  OAI21X1 U3715 ( .A(n4531), .B(n2652), .C(n6400), .Y(n8572) );
  NAND2X1 U3716 ( .A(arr[1814]), .B(n2654), .Y(n6400) );
  OAI21X1 U3718 ( .A(n4467), .B(n2651), .C(n6402), .Y(n8573) );
  NAND2X1 U3719 ( .A(arr[1815]), .B(n2650), .Y(n6402) );
  OAI21X1 U3720 ( .A(n4469), .B(n2649), .C(n6403), .Y(n8574) );
  NAND2X1 U3721 ( .A(arr[1816]), .B(n2650), .Y(n6403) );
  OAI21X1 U3722 ( .A(n4471), .B(n2649), .C(n6404), .Y(n8575) );
  NAND2X1 U3723 ( .A(arr[1817]), .B(n2650), .Y(n6404) );
  OAI21X1 U3724 ( .A(n4473), .B(n2649), .C(n6405), .Y(n8576) );
  NAND2X1 U3725 ( .A(arr[1818]), .B(n2650), .Y(n6405) );
  OAI21X1 U3726 ( .A(n4475), .B(n2649), .C(n6406), .Y(n8577) );
  NAND2X1 U3727 ( .A(arr[1819]), .B(n2650), .Y(n6406) );
  OAI21X1 U3728 ( .A(n4477), .B(n2649), .C(n6407), .Y(n8578) );
  NAND2X1 U3729 ( .A(arr[1820]), .B(n2651), .Y(n6407) );
  OAI21X1 U3730 ( .A(n4479), .B(n2649), .C(n6408), .Y(n8579) );
  NAND2X1 U3731 ( .A(arr[1821]), .B(n2651), .Y(n6408) );
  OAI21X1 U3732 ( .A(n4481), .B(n2650), .C(n6409), .Y(n8580) );
  NAND2X1 U3733 ( .A(arr[1822]), .B(n2650), .Y(n6409) );
  OAI21X1 U3734 ( .A(n4483), .B(n2649), .C(n6410), .Y(n8581) );
  NAND2X1 U3735 ( .A(arr[1823]), .B(n2650), .Y(n6410) );
  OAI21X1 U3736 ( .A(n4485), .B(n2650), .C(n6411), .Y(n8582) );
  NAND2X1 U3737 ( .A(arr[1824]), .B(n2651), .Y(n6411) );
  OAI21X1 U3738 ( .A(n4487), .B(n2650), .C(n6412), .Y(n8583) );
  NAND2X1 U3739 ( .A(arr[1825]), .B(n2651), .Y(n6412) );
  OAI21X1 U3740 ( .A(n4489), .B(n2649), .C(n6413), .Y(n8584) );
  NAND2X1 U3741 ( .A(arr[1826]), .B(n2651), .Y(n6413) );
  OAI21X1 U3742 ( .A(n4491), .B(n2650), .C(n6414), .Y(n8585) );
  NAND2X1 U3743 ( .A(arr[1827]), .B(n2651), .Y(n6414) );
  OAI21X1 U3744 ( .A(n4493), .B(n2650), .C(n6415), .Y(n8586) );
  NAND2X1 U3745 ( .A(arr[1828]), .B(n2651), .Y(n6415) );
  OAI21X1 U3746 ( .A(n4495), .B(n2649), .C(n6416), .Y(n8587) );
  NAND2X1 U3747 ( .A(arr[1829]), .B(n2651), .Y(n6416) );
  OAI21X1 U3748 ( .A(n4497), .B(n2650), .C(n6417), .Y(n8588) );
  NAND2X1 U3749 ( .A(arr[1830]), .B(n2651), .Y(n6417) );
  OAI21X1 U3750 ( .A(n4499), .B(n2650), .C(n6418), .Y(n8589) );
  NAND2X1 U3751 ( .A(arr[1831]), .B(n2651), .Y(n6418) );
  OAI21X1 U3752 ( .A(n4501), .B(n2649), .C(n6419), .Y(n8590) );
  NAND2X1 U3753 ( .A(arr[1832]), .B(n2651), .Y(n6419) );
  OAI21X1 U3754 ( .A(n4503), .B(n2649), .C(n6420), .Y(n8591) );
  NAND2X1 U3755 ( .A(arr[1833]), .B(n2651), .Y(n6420) );
  OAI21X1 U3756 ( .A(n4505), .B(n2649), .C(n6421), .Y(n8592) );
  NAND2X1 U3757 ( .A(arr[1834]), .B(n2651), .Y(n6421) );
  OAI21X1 U3758 ( .A(n4507), .B(n2649), .C(n6422), .Y(n8593) );
  NAND2X1 U3759 ( .A(arr[1835]), .B(n2651), .Y(n6422) );
  OAI21X1 U3760 ( .A(n4509), .B(n2649), .C(n6423), .Y(n8594) );
  NAND2X1 U3761 ( .A(arr[1836]), .B(n2651), .Y(n6423) );
  OAI21X1 U3762 ( .A(n4511), .B(n2649), .C(n6424), .Y(n8595) );
  NAND2X1 U3763 ( .A(arr[1837]), .B(n2651), .Y(n6424) );
  OAI21X1 U3764 ( .A(n4513), .B(n2651), .C(n6425), .Y(n8596) );
  NAND2X1 U3765 ( .A(arr[1838]), .B(n2651), .Y(n6425) );
  OAI21X1 U3766 ( .A(n4515), .B(n2649), .C(n6426), .Y(n8597) );
  NAND2X1 U3767 ( .A(arr[1839]), .B(n2651), .Y(n6426) );
  OAI21X1 U3768 ( .A(n4517), .B(n2650), .C(n6427), .Y(n8598) );
  NAND2X1 U3769 ( .A(arr[1840]), .B(n2651), .Y(n6427) );
  OAI21X1 U3770 ( .A(n4519), .B(n2649), .C(n6428), .Y(n8599) );
  NAND2X1 U3771 ( .A(arr[1841]), .B(n2650), .Y(n6428) );
  OAI21X1 U3772 ( .A(n4521), .B(n2650), .C(n6429), .Y(n8600) );
  NAND2X1 U3773 ( .A(arr[1842]), .B(n2651), .Y(n6429) );
  OAI21X1 U3774 ( .A(n4523), .B(n2649), .C(n6430), .Y(n8601) );
  NAND2X1 U3775 ( .A(arr[1843]), .B(n2650), .Y(n6430) );
  OAI21X1 U3776 ( .A(n4525), .B(n2649), .C(n6431), .Y(n8602) );
  NAND2X1 U3777 ( .A(arr[1844]), .B(n2651), .Y(n6431) );
  OAI21X1 U3778 ( .A(n4527), .B(n2649), .C(n6432), .Y(n8603) );
  NAND2X1 U3779 ( .A(arr[1845]), .B(n2650), .Y(n6432) );
  OAI21X1 U3780 ( .A(n4529), .B(n2649), .C(n6433), .Y(n8604) );
  NAND2X1 U3781 ( .A(arr[1846]), .B(n2650), .Y(n6433) );
  OAI21X1 U3782 ( .A(n4531), .B(n2649), .C(n6434), .Y(n8605) );
  NAND2X1 U3783 ( .A(arr[1847]), .B(n2651), .Y(n6434) );
  AND2X1 U3785 ( .A(n6230), .B(n5887), .Y(n5294) );
  NOR2X1 U3786 ( .A(n6435), .B(wr_ptr[3]), .Y(n6230) );
  AND2X1 U3921 ( .A(n6504), .B(n5680), .Y(n5363) );
  NOR2X1 U3922 ( .A(wr_ptr[1]), .B(wr_ptr[2]), .Y(n5680) );
  AND2X1 U4057 ( .A(n6504), .B(n5749), .Y(n5432) );
  NOR2X1 U4058 ( .A(n6573), .B(wr_ptr[2]), .Y(n5749) );
  AND2X1 U4193 ( .A(n6504), .B(n5818), .Y(n5501) );
  NOR2X1 U4194 ( .A(n6642), .B(wr_ptr[1]), .Y(n5818) );
  AND2X1 U4362 ( .A(n6504), .B(n5887), .Y(n5570) );
  NOR2X1 U4363 ( .A(n6642), .B(n6573), .Y(n5887) );
  NOR2X1 U4364 ( .A(n6435), .B(n6161), .Y(n6504) );
  AND2X1 U4366 ( .A(wr_ptr[5]), .B(n5607), .Y(n6677) );
  OAI21X1 U4368 ( .A(n5608), .B(n6712), .C(n6713), .Y(n8870) );
  NAND2X1 U4369 ( .A(n91), .B(n5607), .Y(n6713) );
  OAI21X1 U4371 ( .A(n6435), .B(n6712), .C(n6714), .Y(n8871) );
  NAND2X1 U4372 ( .A(n90), .B(n5607), .Y(n6714) );
  OAI21X1 U4374 ( .A(n6161), .B(n6712), .C(n6715), .Y(n8872) );
  NAND2X1 U4375 ( .A(n89), .B(n5607), .Y(n6715) );
  OAI21X1 U4377 ( .A(n6642), .B(n6712), .C(n6716), .Y(n8873) );
  NAND2X1 U4378 ( .A(n88), .B(n5607), .Y(n6716) );
  OAI21X1 U4380 ( .A(n6573), .B(n6712), .C(n6717), .Y(n8874) );
  NAND2X1 U4381 ( .A(n87), .B(n5607), .Y(n6717) );
  OAI21X1 U4383 ( .A(n5572), .B(n6712), .C(n6718), .Y(n8875) );
  NAND2X1 U4384 ( .A(n86), .B(n5607), .Y(n6718) );
  NAND2X1 U4386 ( .A(n6719), .B(n6720), .Y(n6712) );
  OAI21X1 U4389 ( .A(n6722), .B(n6723), .C(n6724), .Y(n8876) );
  AOI22X1 U4390 ( .A(n97), .B(n6725), .C(n2224), .D(n6726), .Y(n6724) );
  OAI21X1 U4392 ( .A(n6722), .B(n6727), .C(n6728), .Y(n8877) );
  AOI22X1 U4393 ( .A(n96), .B(n6725), .C(n2223), .D(n6726), .Y(n6728) );
  OAI21X1 U4394 ( .A(n6722), .B(n6729), .C(n6730), .Y(n8878) );
  AOI22X1 U4395 ( .A(n95), .B(n6725), .C(n2222), .D(n6726), .Y(n6730) );
  OAI21X1 U4396 ( .A(n6722), .B(n6731), .C(n6732), .Y(n8879) );
  AOI22X1 U4397 ( .A(n94), .B(n6725), .C(n2221), .D(n6726), .Y(n6732) );
  OAI21X1 U4398 ( .A(n6722), .B(n6733), .C(n6734), .Y(n8880) );
  AOI22X1 U4399 ( .A(n98), .B(n6725), .C(n2225), .D(n6726), .Y(n6734) );
  OAI21X1 U4401 ( .A(n6722), .B(n6735), .C(n6736), .Y(n8881) );
  AOI22X1 U4402 ( .A(n93), .B(n6725), .C(n2220), .D(n6726), .Y(n6736) );
  OAI21X1 U4403 ( .A(n6722), .B(n6737), .C(n6738), .Y(n8882) );
  AOI22X1 U4404 ( .A(n92), .B(n6725), .C(n2219), .D(n6726), .Y(n6738) );
  NAND3X1 U4406 ( .A(n6722), .B(get), .C(n6740), .Y(n6739) );
  NOR2X1 U4407 ( .A(reset), .B(empty), .Y(n6740) );
  NOR2X1 U4408 ( .A(n6741), .B(n4465), .Y(n6725) );
  OAI21X1 U4410 ( .A(n6721), .B(n4465), .C(n6742), .Y(n6741) );
  NAND3X1 U4411 ( .A(n6743), .B(n6720), .C(n6744), .Y(n6742) );
  NOR2X1 U4412 ( .A(n6745), .B(n6746), .Y(n6744) );
  AOI21X1 U4414 ( .A(n6748), .B(n6749), .C(n6750), .Y(n6747) );
  OAI21X1 U4415 ( .A(empty), .B(n6745), .C(n6720), .Y(n4465) );
  NOR2X1 U4418 ( .A(n6746), .B(full), .Y(n6721) );
  NOR2X1 U4420 ( .A(n6749), .B(n6750), .Y(full) );
  NAND3X1 U4421 ( .A(fillcount[1]), .B(n6737), .C(fillcount[2]), .Y(n6749) );
  NOR2X1 U4422 ( .A(n6750), .B(n6748), .Y(empty) );
  NAND3X1 U4423 ( .A(n6735), .B(n6731), .C(n6737), .Y(n6748) );
  NAND3X1 U4427 ( .A(n6729), .B(n6727), .C(n6751), .Y(n6750) );
  NOR2X1 U4428 ( .A(fillcount[6]), .B(fillcount[5]), .Y(n6751) );
  INVX2 U3 ( .A(n4457), .Y(n6752) );
  INVX2 U5 ( .A(n4460), .Y(n6753) );
  INVX2 U7 ( .A(n4461), .Y(n6754) );
  INVX2 U9 ( .A(n4462), .Y(n6755) );
  INVX2 U11 ( .A(n4463), .Y(n6756) );
  INVX2 U13 ( .A(n4464), .Y(n6757) );
  INVX2 U16 ( .A(n4465), .Y(n4459) );
  INVX2 U4265 ( .A(data_in[0]), .Y(n4467) );
  INVX2 U4268 ( .A(data_in[1]), .Y(n4469) );
  INVX2 U4271 ( .A(data_in[2]), .Y(n4471) );
  INVX2 U4274 ( .A(data_in[3]), .Y(n4473) );
  INVX2 U4277 ( .A(data_in[4]), .Y(n4475) );
  INVX2 U4280 ( .A(data_in[5]), .Y(n4477) );
  INVX2 U4283 ( .A(data_in[6]), .Y(n4479) );
  INVX2 U4286 ( .A(data_in[7]), .Y(n4481) );
  INVX2 U4289 ( .A(data_in[8]), .Y(n4483) );
  INVX2 U4292 ( .A(data_in[9]), .Y(n4485) );
  INVX2 U4295 ( .A(data_in[10]), .Y(n4487) );
  INVX2 U4298 ( .A(data_in[11]), .Y(n4489) );
  INVX2 U4301 ( .A(data_in[12]), .Y(n4491) );
  INVX2 U4304 ( .A(data_in[13]), .Y(n4493) );
  INVX2 U4307 ( .A(data_in[14]), .Y(n4495) );
  INVX2 U4310 ( .A(data_in[15]), .Y(n4497) );
  INVX2 U4313 ( .A(data_in[16]), .Y(n4499) );
  INVX2 U4316 ( .A(data_in[17]), .Y(n4501) );
  INVX2 U4319 ( .A(data_in[18]), .Y(n4503) );
  INVX2 U4322 ( .A(data_in[19]), .Y(n4505) );
  INVX2 U4325 ( .A(data_in[20]), .Y(n4507) );
  INVX2 U4328 ( .A(data_in[21]), .Y(n4509) );
  INVX2 U4331 ( .A(data_in[22]), .Y(n4511) );
  INVX2 U4334 ( .A(data_in[23]), .Y(n4513) );
  INVX2 U4337 ( .A(data_in[24]), .Y(n4515) );
  INVX2 U4340 ( .A(data_in[25]), .Y(n4517) );
  INVX2 U4343 ( .A(data_in[26]), .Y(n4519) );
  INVX2 U4346 ( .A(data_in[27]), .Y(n4521) );
  INVX2 U4349 ( .A(data_in[28]), .Y(n4523) );
  INVX2 U4352 ( .A(data_in[29]), .Y(n4525) );
  INVX2 U4355 ( .A(data_in[30]), .Y(n4527) );
  INVX2 U4358 ( .A(data_in[31]), .Y(n4529) );
  INVX2 U4367 ( .A(data_in[32]), .Y(n4531) );
  INVX2 U4370 ( .A(wr_ptr[5]), .Y(n5608) );
  INVX2 U4373 ( .A(wr_ptr[4]), .Y(n6435) );
  INVX2 U4376 ( .A(wr_ptr[3]), .Y(n6161) );
  INVX2 U4379 ( .A(wr_ptr[2]), .Y(n6642) );
  INVX2 U4382 ( .A(wr_ptr[1]), .Y(n6573) );
  INVX2 U4388 ( .A(wr_ptr[0]), .Y(n5572) );
  INVX2 U4400 ( .A(fillcount[6]), .Y(n6733) );
  INVX2 U4405 ( .A(n6739), .Y(n6726) );
  INVX2 U4409 ( .A(n6741), .Y(n6722) );
  INVX2 U4413 ( .A(n6747), .Y(n6743) );
  INVX2 U4416 ( .A(reset), .Y(n6720) );
  INVX2 U4417 ( .A(get), .Y(n6745) );
  INVX2 U4419 ( .A(put), .Y(n6746) );
  INVX2 U4424 ( .A(fillcount[0]), .Y(n6737) );
  INVX2 U4425 ( .A(fillcount[2]), .Y(n6731) );
  INVX2 U4426 ( .A(fillcount[1]), .Y(n6735) );
  INVX2 U4429 ( .A(fillcount[4]), .Y(n6727) );
  INVX2 U4430 ( .A(fillcount[3]), .Y(n6729) );
  FIFO_DEPTH_P26_WIDTH33_DW01_dec_0 sub_55 ( .A(fillcount), .SUM({n2225, n2224, 
        n2223, n2222, n2221, n2220, n2219}) );
  FIFO_DEPTH_P26_WIDTH33_DW01_inc_0 add_54 ( .A({n18, n17, n16, n15, n14, n13}), .SUM({n2218, n2217, n2216, n2215, n2214, n2213}) );
  FIFO_DEPTH_P26_WIDTH33_DW01_inc_1 add_50 ( .A(fillcount), .SUM({n98, n97, 
        n96, n95, n94, n93, n92}) );
  FIFO_DEPTH_P26_WIDTH33_DW01_inc_2 add_49 ( .A(wr_ptr), .SUM({n91, n90, n89, 
        n88, n87, n86}) );
  AND2X2 U83 ( .A(n5570), .B(n4569), .Y(n1) );
  AND2X2 U150 ( .A(n5501), .B(n4569), .Y(n2) );
  AND2X2 U217 ( .A(n5432), .B(n4569), .Y(n3) );
  AND2X2 U284 ( .A(n5363), .B(n4569), .Y(n4) );
  AND2X2 U351 ( .A(n5294), .B(n4569), .Y(n5) );
  AND2X2 U418 ( .A(n5225), .B(n4569), .Y(n6) );
  AND2X2 U485 ( .A(n5156), .B(n4569), .Y(n7) );
  AND2X2 U552 ( .A(n5087), .B(n4569), .Y(n8) );
  AND2X2 U619 ( .A(n5018), .B(n4569), .Y(n9) );
  AND2X2 U686 ( .A(n4949), .B(n4569), .Y(n10) );
  AND2X2 U753 ( .A(n4880), .B(n4569), .Y(n11) );
  AND2X2 U820 ( .A(n4811), .B(n4569), .Y(n12) );
  AND2X2 U887 ( .A(n4742), .B(n4569), .Y(n19) );
  AND2X2 U954 ( .A(n4673), .B(n4569), .Y(n20) );
  AND2X2 U1021 ( .A(n4604), .B(n4569), .Y(n21) );
  AND2X2 U1088 ( .A(n4569), .B(n4534), .Y(n22) );
  AND2X2 U1155 ( .A(n5678), .B(n5294), .Y(n23) );
  AND2X2 U1222 ( .A(n5678), .B(n5225), .Y(n24) );
  AND2X2 U1289 ( .A(n5678), .B(n5156), .Y(n25) );
  AND2X2 U1356 ( .A(n5678), .B(n5087), .Y(n26) );
  AND2X2 U1423 ( .A(n5678), .B(n5018), .Y(n27) );
  AND2X2 U1490 ( .A(n5678), .B(n4949), .Y(n28) );
  AND2X2 U1557 ( .A(n5678), .B(n4880), .Y(n29) );
  AND2X2 U1624 ( .A(n5678), .B(n4811), .Y(n30) );
  AND2X2 U1691 ( .A(n5678), .B(n4742), .Y(n31) );
  AND2X2 U1758 ( .A(n5678), .B(n4673), .Y(n32) );
  AND2X2 U1825 ( .A(n5678), .B(n4604), .Y(n33) );
  AND2X2 U1892 ( .A(n5678), .B(n4534), .Y(n34) );
  AND2X2 U1959 ( .A(n5643), .B(n5294), .Y(n35) );
  AND2X2 U2026 ( .A(n5643), .B(n5225), .Y(n36) );
  AND2X2 U2093 ( .A(n5643), .B(n5156), .Y(n37) );
  AND2X2 U2094 ( .A(n5643), .B(n5087), .Y(n38) );
  AND2X2 U2161 ( .A(n5643), .B(n5018), .Y(n39) );
  AND2X2 U2162 ( .A(n5643), .B(n4949), .Y(n40) );
  AND2X2 U2230 ( .A(n5643), .B(n4880), .Y(n41) );
  AND2X2 U2297 ( .A(n5643), .B(n4811), .Y(n42) );
  AND2X2 U2365 ( .A(n5643), .B(n4742), .Y(n43) );
  AND2X2 U2432 ( .A(n5643), .B(n4673), .Y(n44) );
  AND2X2 U2500 ( .A(n5643), .B(n4604), .Y(n45) );
  AND2X2 U2567 ( .A(n5643), .B(n4534), .Y(n46) );
  INVX2 U2635 ( .A(n22), .Y(n2813) );
  INVX2 U2702 ( .A(n22), .Y(n2812) );
  INVX2 U2771 ( .A(n23), .Y(n2651) );
  INVX2 U2838 ( .A(n23), .Y(n2650) );
  INVX2 U2906 ( .A(n35), .Y(n2654) );
  INVX2 U2973 ( .A(n35), .Y(n2653) );
  INVX2 U3041 ( .A(n24), .Y(n2657) );
  INVX2 U3108 ( .A(n24), .Y(n2656) );
  INVX2 U3176 ( .A(n36), .Y(n2660) );
  INVX2 U3243 ( .A(n36), .Y(n2659) );
  INVX2 U3312 ( .A(n25), .Y(n2663) );
  INVX2 U3379 ( .A(n25), .Y(n2662) );
  INVX2 U3447 ( .A(n37), .Y(n2666) );
  INVX2 U3514 ( .A(n37), .Y(n2665) );
  INVX2 U3582 ( .A(n26), .Y(n2669) );
  INVX2 U3649 ( .A(n26), .Y(n2668) );
  INVX2 U3717 ( .A(n38), .Y(n2672) );
  INVX2 U3784 ( .A(n38), .Y(n2671) );
  INVX2 U3787 ( .A(n27), .Y(n2675) );
  INVX2 U3788 ( .A(n27), .Y(n2674) );
  INVX2 U3789 ( .A(n39), .Y(n2678) );
  INVX2 U3790 ( .A(n39), .Y(n2677) );
  INVX2 U3791 ( .A(n28), .Y(n2681) );
  INVX2 U3792 ( .A(n28), .Y(n2680) );
  INVX2 U3793 ( .A(n40), .Y(n2684) );
  INVX2 U3794 ( .A(n40), .Y(n2683) );
  INVX2 U3795 ( .A(n29), .Y(n2687) );
  INVX2 U3796 ( .A(n29), .Y(n2686) );
  INVX2 U3797 ( .A(n41), .Y(n2690) );
  INVX2 U3798 ( .A(n41), .Y(n2689) );
  INVX2 U3799 ( .A(n30), .Y(n2693) );
  INVX2 U3800 ( .A(n30), .Y(n2692) );
  INVX2 U3801 ( .A(n42), .Y(n2696) );
  INVX2 U3802 ( .A(n42), .Y(n2695) );
  INVX2 U3803 ( .A(n31), .Y(n2699) );
  INVX2 U3804 ( .A(n31), .Y(n2698) );
  INVX2 U3805 ( .A(n43), .Y(n2702) );
  INVX2 U3806 ( .A(n43), .Y(n2701) );
  INVX2 U3807 ( .A(n32), .Y(n2705) );
  INVX2 U3808 ( .A(n32), .Y(n2704) );
  INVX2 U3809 ( .A(n44), .Y(n2708) );
  INVX2 U3810 ( .A(n44), .Y(n2707) );
  INVX2 U3811 ( .A(n33), .Y(n2711) );
  INVX2 U3812 ( .A(n33), .Y(n2710) );
  INVX2 U3813 ( .A(n45), .Y(n2714) );
  INVX2 U3814 ( .A(n45), .Y(n2713) );
  INVX2 U3815 ( .A(n34), .Y(n2717) );
  INVX2 U3816 ( .A(n34), .Y(n2716) );
  INVX2 U3817 ( .A(n46), .Y(n2720) );
  INVX2 U3818 ( .A(n46), .Y(n2719) );
  INVX2 U3819 ( .A(n1), .Y(n2723) );
  INVX2 U3820 ( .A(n1), .Y(n2722) );
  INVX2 U3821 ( .A(n2), .Y(n2729) );
  INVX2 U3822 ( .A(n2), .Y(n2728) );
  INVX2 U3823 ( .A(n3), .Y(n2735) );
  INVX2 U3824 ( .A(n3), .Y(n2734) );
  INVX2 U3825 ( .A(n4), .Y(n2741) );
  INVX2 U3826 ( .A(n4), .Y(n2740) );
  INVX2 U3827 ( .A(n5), .Y(n2747) );
  INVX2 U3828 ( .A(n5), .Y(n2746) );
  INVX2 U3829 ( .A(n6), .Y(n2753) );
  INVX2 U3830 ( .A(n6), .Y(n2752) );
  INVX2 U3831 ( .A(n7), .Y(n2759) );
  INVX2 U3832 ( .A(n7), .Y(n2758) );
  INVX2 U3833 ( .A(n8), .Y(n2765) );
  INVX2 U3834 ( .A(n8), .Y(n2764) );
  INVX2 U3835 ( .A(n9), .Y(n2771) );
  INVX2 U3836 ( .A(n9), .Y(n2770) );
  INVX2 U3837 ( .A(n10), .Y(n2777) );
  INVX2 U3838 ( .A(n10), .Y(n2776) );
  INVX2 U3839 ( .A(n11), .Y(n2783) );
  INVX2 U3840 ( .A(n11), .Y(n2782) );
  INVX2 U3841 ( .A(n12), .Y(n2789) );
  INVX2 U3842 ( .A(n12), .Y(n2788) );
  INVX2 U3843 ( .A(n19), .Y(n2795) );
  INVX2 U3844 ( .A(n19), .Y(n2794) );
  INVX2 U3845 ( .A(n20), .Y(n2801) );
  INVX2 U3846 ( .A(n20), .Y(n2800) );
  INVX2 U3847 ( .A(n21), .Y(n2807) );
  INVX2 U3848 ( .A(n21), .Y(n2806) );
  AND2X2 U3849 ( .A(n5570), .B(n4533), .Y(n47) );
  AND2X2 U3850 ( .A(n5501), .B(n4533), .Y(n48) );
  AND2X2 U3851 ( .A(n5432), .B(n4533), .Y(n49) );
  AND2X2 U3852 ( .A(n5363), .B(n4533), .Y(n50) );
  AND2X2 U3853 ( .A(n5294), .B(n4533), .Y(n51) );
  AND2X2 U3854 ( .A(n5225), .B(n4533), .Y(n52) );
  AND2X2 U3855 ( .A(n5156), .B(n4533), .Y(n53) );
  AND2X2 U3856 ( .A(n5087), .B(n4533), .Y(n54) );
  AND2X2 U3857 ( .A(n5018), .B(n4533), .Y(n55) );
  AND2X2 U3858 ( .A(n4949), .B(n4533), .Y(n56) );
  AND2X2 U3859 ( .A(n4880), .B(n4533), .Y(n57) );
  AND2X2 U3860 ( .A(n4811), .B(n4533), .Y(n58) );
  AND2X2 U3861 ( .A(n4742), .B(n4533), .Y(n59) );
  AND2X2 U3862 ( .A(n4673), .B(n4533), .Y(n60) );
  AND2X2 U3863 ( .A(n4604), .B(n4533), .Y(n61) );
  AND2X2 U3864 ( .A(n4533), .B(n4534), .Y(n62) );
  AND2X2 U3865 ( .A(n5643), .B(n5363), .Y(n63) );
  AND2X2 U3866 ( .A(n5678), .B(n5363), .Y(n64) );
  AND2X2 U3867 ( .A(n5643), .B(n5432), .Y(n65) );
  AND2X2 U3868 ( .A(n5678), .B(n5432), .Y(n66) );
  AND2X2 U3869 ( .A(n5643), .B(n5501), .Y(n67) );
  AND2X2 U3870 ( .A(n5678), .B(n5501), .Y(n68) );
  AND2X2 U3871 ( .A(n5643), .B(n5570), .Y(n69) );
  AND2X2 U3872 ( .A(n5678), .B(n5570), .Y(n70) );
  INVX2 U3873 ( .A(n46), .Y(n2718) );
  INVX2 U3874 ( .A(n45), .Y(n2712) );
  INVX2 U3875 ( .A(n44), .Y(n2706) );
  INVX2 U3876 ( .A(n43), .Y(n2700) );
  INVX2 U3877 ( .A(n42), .Y(n2694) );
  INVX2 U3878 ( .A(n41), .Y(n2688) );
  INVX2 U3879 ( .A(n40), .Y(n2682) );
  INVX2 U3880 ( .A(n39), .Y(n2676) );
  INVX2 U3881 ( .A(n38), .Y(n2670) );
  INVX2 U3882 ( .A(n37), .Y(n2664) );
  INVX2 U3883 ( .A(n36), .Y(n2658) );
  INVX2 U3884 ( .A(n35), .Y(n2652) );
  INVX2 U3885 ( .A(n61), .Y(n2809) );
  INVX2 U3886 ( .A(n61), .Y(n2808) );
  INVX2 U3887 ( .A(n60), .Y(n2803) );
  INVX2 U3888 ( .A(n60), .Y(n2802) );
  INVX2 U3889 ( .A(n59), .Y(n2797) );
  INVX2 U3890 ( .A(n59), .Y(n2796) );
  INVX2 U3891 ( .A(n58), .Y(n2791) );
  INVX2 U3892 ( .A(n58), .Y(n2790) );
  INVX2 U3893 ( .A(n57), .Y(n2785) );
  INVX2 U3894 ( .A(n57), .Y(n2784) );
  INVX2 U3895 ( .A(n56), .Y(n2779) );
  INVX2 U3896 ( .A(n56), .Y(n2778) );
  INVX2 U3897 ( .A(n55), .Y(n2773) );
  INVX2 U3898 ( .A(n55), .Y(n2772) );
  INVX2 U3899 ( .A(n54), .Y(n2767) );
  INVX2 U3900 ( .A(n54), .Y(n2766) );
  INVX2 U3901 ( .A(n53), .Y(n2761) );
  INVX2 U3902 ( .A(n53), .Y(n2760) );
  INVX2 U3903 ( .A(n52), .Y(n2755) );
  INVX2 U3904 ( .A(n52), .Y(n2754) );
  INVX2 U3905 ( .A(n51), .Y(n2749) );
  INVX2 U3906 ( .A(n51), .Y(n2748) );
  INVX2 U3907 ( .A(n50), .Y(n2743) );
  INVX2 U3908 ( .A(n50), .Y(n2742) );
  INVX2 U3909 ( .A(n49), .Y(n2737) );
  INVX2 U3910 ( .A(n49), .Y(n2736) );
  INVX2 U3911 ( .A(n48), .Y(n2731) );
  INVX2 U3912 ( .A(n48), .Y(n2730) );
  INVX2 U3913 ( .A(n47), .Y(n2725) );
  INVX2 U3914 ( .A(n47), .Y(n2724) );
  INVX2 U3915 ( .A(n61), .Y(n2810) );
  INVX2 U3916 ( .A(n60), .Y(n2804) );
  INVX2 U3917 ( .A(n59), .Y(n2798) );
  INVX2 U3918 ( .A(n58), .Y(n2792) );
  INVX2 U3919 ( .A(n57), .Y(n2786) );
  INVX2 U3920 ( .A(n56), .Y(n2780) );
  INVX2 U3923 ( .A(n55), .Y(n2774) );
  INVX2 U3924 ( .A(n54), .Y(n2768) );
  INVX2 U3925 ( .A(n53), .Y(n2762) );
  INVX2 U3926 ( .A(n52), .Y(n2756) );
  INVX2 U3927 ( .A(n51), .Y(n2750) );
  INVX2 U3928 ( .A(n50), .Y(n2744) );
  INVX2 U3929 ( .A(n49), .Y(n2738) );
  INVX2 U3930 ( .A(n48), .Y(n2732) );
  INVX2 U3931 ( .A(n47), .Y(n2726) );
  INVX2 U3932 ( .A(n62), .Y(n2815) );
  INVX2 U3933 ( .A(n62), .Y(n2814) );
  INVX2 U3934 ( .A(n62), .Y(n2816) );
  INVX2 U3935 ( .A(n22), .Y(n2811) );
  INVX2 U3936 ( .A(n34), .Y(n2715) );
  INVX2 U3937 ( .A(n33), .Y(n2709) );
  INVX2 U3938 ( .A(n32), .Y(n2703) );
  INVX2 U3939 ( .A(n31), .Y(n2697) );
  INVX2 U3940 ( .A(n30), .Y(n2691) );
  INVX2 U3941 ( .A(n29), .Y(n2685) );
  INVX2 U3942 ( .A(n28), .Y(n2679) );
  INVX2 U3943 ( .A(n27), .Y(n2673) );
  INVX2 U3944 ( .A(n26), .Y(n2667) );
  INVX2 U3945 ( .A(n25), .Y(n2661) );
  INVX2 U3946 ( .A(n24), .Y(n2655) );
  INVX2 U3947 ( .A(n23), .Y(n2649) );
  INVX2 U3948 ( .A(n21), .Y(n2805) );
  INVX2 U3949 ( .A(n20), .Y(n2799) );
  INVX2 U3950 ( .A(n19), .Y(n2793) );
  INVX2 U3951 ( .A(n12), .Y(n2787) );
  INVX2 U3952 ( .A(n11), .Y(n2781) );
  INVX2 U3953 ( .A(n10), .Y(n2775) );
  INVX2 U3954 ( .A(n9), .Y(n2769) );
  INVX2 U3955 ( .A(n8), .Y(n2763) );
  INVX2 U3956 ( .A(n7), .Y(n2757) );
  INVX2 U3957 ( .A(n6), .Y(n2751) );
  INVX2 U3958 ( .A(n5), .Y(n2745) );
  INVX2 U3959 ( .A(n4), .Y(n2739) );
  INVX2 U3960 ( .A(n3), .Y(n2733) );
  INVX2 U3961 ( .A(n2), .Y(n2727) );
  INVX2 U3962 ( .A(n1), .Y(n2721) );
  INVX2 U3963 ( .A(n63), .Y(n2648) );
  INVX2 U3964 ( .A(n65), .Y(n2646) );
  INVX2 U3965 ( .A(n67), .Y(n2644) );
  INVX2 U3966 ( .A(n69), .Y(n2642) );
  BUFX2 U3967 ( .A(n2436), .Y(n2437) );
  BUFX2 U3968 ( .A(n2436), .Y(n2438) );
  BUFX2 U3969 ( .A(n2435), .Y(n2440) );
  BUFX2 U3970 ( .A(n2436), .Y(n2439) );
  BUFX2 U3971 ( .A(n2435), .Y(n2441) );
  BUFX2 U3972 ( .A(n2435), .Y(n2442) );
  BUFX2 U3973 ( .A(n2434), .Y(n2444) );
  BUFX2 U3974 ( .A(n2434), .Y(n2443) );
  BUFX2 U3975 ( .A(n2434), .Y(n2445) );
  BUFX2 U3976 ( .A(n2433), .Y(n2446) );
  BUFX2 U3977 ( .A(n2433), .Y(n2448) );
  BUFX2 U3978 ( .A(n2433), .Y(n2447) );
  BUFX2 U3979 ( .A(n2432), .Y(n2449) );
  BUFX2 U3980 ( .A(n2432), .Y(n2450) );
  BUFX2 U3981 ( .A(n2431), .Y(n2452) );
  BUFX2 U3982 ( .A(n2432), .Y(n2451) );
  BUFX2 U3983 ( .A(n2431), .Y(n2453) );
  BUFX2 U3984 ( .A(n2431), .Y(n2454) );
  BUFX2 U3985 ( .A(n2430), .Y(n2456) );
  BUFX2 U3986 ( .A(n2430), .Y(n2455) );
  BUFX2 U3987 ( .A(n2430), .Y(n2457) );
  BUFX2 U3988 ( .A(n2429), .Y(n2458) );
  BUFX2 U3989 ( .A(n2429), .Y(n2460) );
  BUFX2 U3990 ( .A(n2429), .Y(n2459) );
  BUFX2 U3991 ( .A(n2428), .Y(n2461) );
  BUFX2 U3992 ( .A(n2428), .Y(n2462) );
  BUFX2 U3993 ( .A(n2427), .Y(n2464) );
  BUFX2 U3994 ( .A(n2428), .Y(n2463) );
  BUFX2 U3995 ( .A(n2427), .Y(n2465) );
  BUFX2 U3996 ( .A(n2427), .Y(n2466) );
  BUFX2 U3997 ( .A(n2426), .Y(n2468) );
  BUFX2 U3998 ( .A(n2426), .Y(n2467) );
  BUFX2 U3999 ( .A(n2426), .Y(n2469) );
  BUFX2 U4000 ( .A(n2425), .Y(n2470) );
  BUFX2 U4001 ( .A(n2425), .Y(n2472) );
  BUFX2 U4002 ( .A(n2425), .Y(n2471) );
  BUFX2 U4003 ( .A(n2424), .Y(n2473) );
  BUFX2 U4004 ( .A(n2424), .Y(n2474) );
  BUFX2 U4005 ( .A(n2423), .Y(n2476) );
  BUFX2 U4006 ( .A(n2424), .Y(n2475) );
  BUFX2 U4007 ( .A(n2423), .Y(n2477) );
  BUFX2 U4008 ( .A(n2423), .Y(n2478) );
  BUFX2 U4009 ( .A(n2422), .Y(n2480) );
  BUFX2 U4010 ( .A(n2422), .Y(n2479) );
  BUFX2 U4011 ( .A(n2422), .Y(n2481) );
  BUFX2 U4012 ( .A(n2421), .Y(n2482) );
  BUFX2 U4013 ( .A(n2421), .Y(n2484) );
  BUFX2 U4014 ( .A(n2421), .Y(n2483) );
  BUFX2 U4015 ( .A(n2420), .Y(n2485) );
  BUFX2 U4016 ( .A(n2420), .Y(n2486) );
  BUFX2 U4017 ( .A(n2419), .Y(n2488) );
  BUFX2 U4018 ( .A(n2420), .Y(n2487) );
  BUFX2 U4019 ( .A(n2419), .Y(n2489) );
  BUFX2 U4020 ( .A(n2419), .Y(n2490) );
  BUFX2 U4021 ( .A(n2418), .Y(n2492) );
  BUFX2 U4022 ( .A(n2418), .Y(n2491) );
  BUFX2 U4023 ( .A(n2418), .Y(n2493) );
  BUFX2 U4024 ( .A(n2417), .Y(n2494) );
  BUFX2 U4025 ( .A(n2417), .Y(n2496) );
  BUFX2 U4026 ( .A(n2417), .Y(n2495) );
  BUFX2 U4027 ( .A(n2416), .Y(n2497) );
  BUFX2 U4028 ( .A(n2416), .Y(n2498) );
  BUFX2 U4029 ( .A(n2415), .Y(n2500) );
  BUFX2 U4030 ( .A(n2416), .Y(n2499) );
  BUFX2 U4031 ( .A(n2415), .Y(n2501) );
  BUFX2 U4032 ( .A(n2415), .Y(n2502) );
  BUFX2 U4033 ( .A(n2414), .Y(n2504) );
  BUFX2 U4034 ( .A(n2414), .Y(n2503) );
  BUFX2 U4035 ( .A(n2414), .Y(n2505) );
  BUFX2 U4036 ( .A(n2413), .Y(n2506) );
  BUFX2 U4037 ( .A(n2413), .Y(n2508) );
  BUFX2 U4038 ( .A(n2413), .Y(n2507) );
  BUFX2 U4039 ( .A(n2412), .Y(n2509) );
  BUFX2 U4040 ( .A(n2412), .Y(n2510) );
  BUFX2 U4041 ( .A(n2411), .Y(n2512) );
  BUFX2 U4042 ( .A(n2412), .Y(n2511) );
  BUFX2 U4043 ( .A(n2411), .Y(n2513) );
  BUFX2 U4044 ( .A(n2411), .Y(n2514) );
  BUFX2 U4045 ( .A(n2410), .Y(n2516) );
  BUFX2 U4046 ( .A(n2410), .Y(n2515) );
  BUFX2 U4047 ( .A(n2410), .Y(n2517) );
  BUFX2 U4048 ( .A(n2409), .Y(n2518) );
  BUFX2 U4049 ( .A(n2409), .Y(n2520) );
  BUFX2 U4050 ( .A(n2409), .Y(n2519) );
  BUFX2 U4051 ( .A(n2408), .Y(n2521) );
  BUFX2 U4052 ( .A(n2408), .Y(n2522) );
  BUFX2 U4053 ( .A(n2408), .Y(n2523) );
  INVX2 U4054 ( .A(n64), .Y(n2647) );
  INVX2 U4055 ( .A(n66), .Y(n2645) );
  INVX2 U4056 ( .A(n68), .Y(n2643) );
  INVX2 U4059 ( .A(n70), .Y(n2641) );
  BUFX2 U4060 ( .A(n2407), .Y(n2524) );
  BUFX2 U4061 ( .A(n2525), .Y(n2407) );
  BUFX2 U4062 ( .A(n2579), .Y(n2535) );
  BUFX2 U4063 ( .A(n2579), .Y(n2536) );
  BUFX2 U4064 ( .A(n2580), .Y(n2537) );
  BUFX2 U4065 ( .A(n2580), .Y(n2538) );
  BUFX2 U4066 ( .A(n2580), .Y(n2539) );
  BUFX2 U4067 ( .A(n2581), .Y(n2540) );
  BUFX2 U4068 ( .A(n2581), .Y(n2541) );
  BUFX2 U4069 ( .A(n2581), .Y(n2542) );
  BUFX2 U4070 ( .A(n2582), .Y(n2543) );
  BUFX2 U4071 ( .A(n2582), .Y(n2544) );
  BUFX2 U4072 ( .A(n2582), .Y(n2545) );
  BUFX2 U4073 ( .A(n2583), .Y(n2546) );
  BUFX2 U4074 ( .A(n2583), .Y(n2547) );
  BUFX2 U4075 ( .A(n2583), .Y(n2548) );
  BUFX2 U4076 ( .A(n2584), .Y(n2549) );
  BUFX2 U4077 ( .A(n2584), .Y(n2550) );
  BUFX2 U4078 ( .A(n2584), .Y(n2551) );
  BUFX2 U4079 ( .A(n2585), .Y(n2552) );
  BUFX2 U4080 ( .A(n2585), .Y(n2553) );
  BUFX2 U4081 ( .A(n2585), .Y(n2554) );
  BUFX2 U4082 ( .A(n2586), .Y(n2555) );
  BUFX2 U4083 ( .A(n2586), .Y(n2556) );
  BUFX2 U4084 ( .A(n2586), .Y(n2557) );
  BUFX2 U4085 ( .A(n2587), .Y(n2558) );
  BUFX2 U4086 ( .A(n2587), .Y(n2559) );
  BUFX2 U4087 ( .A(n2587), .Y(n2560) );
  BUFX2 U4088 ( .A(n2588), .Y(n2561) );
  BUFX2 U4089 ( .A(n2588), .Y(n2562) );
  BUFX2 U4090 ( .A(n2588), .Y(n2563) );
  BUFX2 U4091 ( .A(n2589), .Y(n2564) );
  BUFX2 U4092 ( .A(n2589), .Y(n2565) );
  BUFX2 U4093 ( .A(n2589), .Y(n2566) );
  BUFX2 U4094 ( .A(n2590), .Y(n2567) );
  BUFX2 U4095 ( .A(n2590), .Y(n2568) );
  BUFX2 U4096 ( .A(n2590), .Y(n2569) );
  BUFX2 U4097 ( .A(n2591), .Y(n2570) );
  BUFX2 U4098 ( .A(n2591), .Y(n2571) );
  BUFX2 U4099 ( .A(n2591), .Y(n2572) );
  BUFX2 U4100 ( .A(n2592), .Y(n2573) );
  BUFX2 U4101 ( .A(n2592), .Y(n2574) );
  BUFX2 U4102 ( .A(n2592), .Y(n2575) );
  BUFX2 U4103 ( .A(n2593), .Y(n2576) );
  BUFX2 U4104 ( .A(n2593), .Y(n2577) );
  BUFX2 U4105 ( .A(n2593), .Y(n2578) );
  BUFX2 U4106 ( .A(n2534), .Y(n2436) );
  BUFX2 U4107 ( .A(n2534), .Y(n2435) );
  BUFX2 U4108 ( .A(n2534), .Y(n2434) );
  BUFX2 U4109 ( .A(n2533), .Y(n2433) );
  BUFX2 U4110 ( .A(n2533), .Y(n2432) );
  BUFX2 U4111 ( .A(n2533), .Y(n2431) );
  BUFX2 U4112 ( .A(n2532), .Y(n2430) );
  BUFX2 U4113 ( .A(n2532), .Y(n2429) );
  BUFX2 U4114 ( .A(n2532), .Y(n2428) );
  BUFX2 U4115 ( .A(n2531), .Y(n2427) );
  BUFX2 U4116 ( .A(n2531), .Y(n2426) );
  BUFX2 U4117 ( .A(n2531), .Y(n2425) );
  BUFX2 U4118 ( .A(n2530), .Y(n2424) );
  BUFX2 U4119 ( .A(n2530), .Y(n2423) );
  BUFX2 U4120 ( .A(n2530), .Y(n2422) );
  BUFX2 U4121 ( .A(n2529), .Y(n2421) );
  BUFX2 U4122 ( .A(n2529), .Y(n2420) );
  BUFX2 U4123 ( .A(n2529), .Y(n2419) );
  BUFX2 U4124 ( .A(n2528), .Y(n2418) );
  BUFX2 U4125 ( .A(n2528), .Y(n2417) );
  BUFX2 U4126 ( .A(n2528), .Y(n2416) );
  BUFX2 U4127 ( .A(n2527), .Y(n2415) );
  BUFX2 U4128 ( .A(n2527), .Y(n2414) );
  BUFX2 U4129 ( .A(n2527), .Y(n2413) );
  BUFX2 U4130 ( .A(n2526), .Y(n2412) );
  BUFX2 U4131 ( .A(n2526), .Y(n2411) );
  BUFX2 U4132 ( .A(n2526), .Y(n2410) );
  BUFX2 U4133 ( .A(n2525), .Y(n2409) );
  BUFX2 U4134 ( .A(n2525), .Y(n2408) );
  BUFX2 U4135 ( .A(n2617), .Y(n2595) );
  BUFX2 U4136 ( .A(n2617), .Y(n2596) );
  BUFX2 U4137 ( .A(n2617), .Y(n2597) );
  BUFX2 U4138 ( .A(n2618), .Y(n2598) );
  BUFX2 U4139 ( .A(n2618), .Y(n2599) );
  BUFX2 U4140 ( .A(n2618), .Y(n2600) );
  BUFX2 U4141 ( .A(n2619), .Y(n2601) );
  BUFX2 U4142 ( .A(n2619), .Y(n2602) );
  BUFX2 U4143 ( .A(n2619), .Y(n2603) );
  BUFX2 U4144 ( .A(n2620), .Y(n2604) );
  BUFX2 U4145 ( .A(n2620), .Y(n2605) );
  BUFX2 U4146 ( .A(n2620), .Y(n2606) );
  BUFX2 U4147 ( .A(n2621), .Y(n2607) );
  BUFX2 U4148 ( .A(n2621), .Y(n2608) );
  BUFX2 U4149 ( .A(n2621), .Y(n2609) );
  BUFX2 U4150 ( .A(n2622), .Y(n2610) );
  BUFX2 U4151 ( .A(n2622), .Y(n2611) );
  BUFX2 U4152 ( .A(n2622), .Y(n2612) );
  BUFX2 U4153 ( .A(n2623), .Y(n2613) );
  BUFX2 U4154 ( .A(n2623), .Y(n2614) );
  BUFX2 U4155 ( .A(n2623), .Y(n2615) );
  BUFX2 U4156 ( .A(n16), .Y(n2624) );
  BUFX2 U4157 ( .A(n16), .Y(n2625) );
  BUFX2 U4158 ( .A(n16), .Y(n2626) );
  BUFX2 U4159 ( .A(n16), .Y(n2627) );
  BUFX2 U4160 ( .A(n16), .Y(n2628) );
  BUFX2 U4161 ( .A(n16), .Y(n2629) );
  BUFX2 U4162 ( .A(n16), .Y(n2630) );
  BUFX2 U4163 ( .A(n16), .Y(n2631) );
  BUFX2 U4164 ( .A(n16), .Y(n2632) );
  BUFX2 U4165 ( .A(n16), .Y(n2633) );
  BUFX2 U4166 ( .A(n16), .Y(n2634) );
  BUFX2 U4167 ( .A(n14), .Y(n2580) );
  BUFX2 U4168 ( .A(n14), .Y(n2581) );
  BUFX2 U4169 ( .A(n14), .Y(n2582) );
  BUFX2 U4170 ( .A(n14), .Y(n2583) );
  BUFX2 U4171 ( .A(n14), .Y(n2584) );
  BUFX2 U4172 ( .A(n14), .Y(n2585) );
  BUFX2 U4173 ( .A(n14), .Y(n2586) );
  BUFX2 U4174 ( .A(n14), .Y(n2587) );
  BUFX2 U4175 ( .A(n14), .Y(n2588) );
  BUFX2 U4176 ( .A(n14), .Y(n2589) );
  BUFX2 U4177 ( .A(n14), .Y(n2590) );
  BUFX2 U4178 ( .A(n14), .Y(n2591) );
  BUFX2 U4179 ( .A(n14), .Y(n2592) );
  BUFX2 U4180 ( .A(n14), .Y(n2593) );
  BUFX2 U4181 ( .A(n13), .Y(n2534) );
  BUFX2 U4182 ( .A(n13), .Y(n2533) );
  BUFX2 U4183 ( .A(n13), .Y(n2532) );
  BUFX2 U4184 ( .A(n13), .Y(n2531) );
  BUFX2 U4185 ( .A(n13), .Y(n2530) );
  BUFX2 U4186 ( .A(n13), .Y(n2529) );
  BUFX2 U4187 ( .A(n13), .Y(n2528) );
  BUFX2 U4188 ( .A(n13), .Y(n2527) );
  BUFX2 U4189 ( .A(n13), .Y(n2526) );
  BUFX2 U4190 ( .A(n13), .Y(n2525) );
  BUFX2 U4191 ( .A(n14), .Y(n2579) );
  AND2X1 U4192 ( .A(arr[1853]), .B(n2648), .Y(n71) );
  AND2X1 U4195 ( .A(arr[1854]), .B(n2648), .Y(n72) );
  AND2X1 U4196 ( .A(arr[1857]), .B(n2648), .Y(n73) );
  AND2X1 U4197 ( .A(arr[1858]), .B(n2648), .Y(n74) );
  AND2X1 U4198 ( .A(arr[1859]), .B(n2648), .Y(n75) );
  AND2X1 U4199 ( .A(arr[1860]), .B(n2648), .Y(n76) );
  AND2X1 U4200 ( .A(arr[1861]), .B(n2648), .Y(n77) );
  AND2X1 U4201 ( .A(arr[1862]), .B(n2648), .Y(n78) );
  AND2X1 U4202 ( .A(arr[1863]), .B(n2648), .Y(n79) );
  AND2X1 U4203 ( .A(arr[1864]), .B(n2648), .Y(n80) );
  AND2X1 U4204 ( .A(arr[1865]), .B(n2648), .Y(n81) );
  AND2X1 U4205 ( .A(arr[1866]), .B(n2648), .Y(n82) );
  AND2X1 U4206 ( .A(arr[1867]), .B(n2648), .Y(n83) );
  AND2X1 U4207 ( .A(arr[1868]), .B(n2648), .Y(n84) );
  AND2X1 U4208 ( .A(arr[1869]), .B(n2648), .Y(n85) );
  AND2X1 U4209 ( .A(arr[1870]), .B(n2648), .Y(n99) );
  AND2X1 U4210 ( .A(arr[1880]), .B(n2648), .Y(n100) );
  AND2X1 U4211 ( .A(arr[1886]), .B(n2647), .Y(n101) );
  AND2X1 U4212 ( .A(arr[1887]), .B(n2647), .Y(n102) );
  AND2X1 U4213 ( .A(arr[1890]), .B(n2647), .Y(n103) );
  AND2X1 U4214 ( .A(arr[1891]), .B(n2647), .Y(n104) );
  AND2X1 U4215 ( .A(arr[1892]), .B(n2647), .Y(n105) );
  AND2X1 U4216 ( .A(arr[1893]), .B(n2647), .Y(n106) );
  AND2X1 U4217 ( .A(arr[1894]), .B(n2647), .Y(n107) );
  AND2X1 U4218 ( .A(arr[1895]), .B(n2647), .Y(n108) );
  AND2X1 U4219 ( .A(arr[1896]), .B(n2647), .Y(n109) );
  AND2X1 U4220 ( .A(arr[1897]), .B(n2647), .Y(n110) );
  AND2X1 U4221 ( .A(arr[1898]), .B(n2647), .Y(n111) );
  AND2X1 U4222 ( .A(arr[1899]), .B(n2647), .Y(n112) );
  AND2X1 U4223 ( .A(arr[1900]), .B(n2647), .Y(n113) );
  AND2X1 U4224 ( .A(arr[1901]), .B(n2647), .Y(n114) );
  AND2X1 U4225 ( .A(arr[1902]), .B(n2647), .Y(n115) );
  AND2X1 U4226 ( .A(arr[1903]), .B(n2647), .Y(n116) );
  AND2X1 U4227 ( .A(arr[1913]), .B(n2647), .Y(n117) );
  AND2X1 U4228 ( .A(arr[1919]), .B(n2646), .Y(n118) );
  AND2X1 U4229 ( .A(arr[1920]), .B(n2646), .Y(n119) );
  AND2X1 U4230 ( .A(arr[1923]), .B(n2646), .Y(n120) );
  AND2X1 U4231 ( .A(arr[1924]), .B(n2646), .Y(n121) );
  AND2X1 U4232 ( .A(arr[1925]), .B(n2646), .Y(n122) );
  AND2X1 U4233 ( .A(arr[1926]), .B(n2646), .Y(n123) );
  AND2X1 U4234 ( .A(arr[1927]), .B(n2646), .Y(n124) );
  AND2X1 U4235 ( .A(arr[1928]), .B(n2646), .Y(n125) );
  AND2X1 U4236 ( .A(arr[1929]), .B(n2646), .Y(n126) );
  AND2X1 U4237 ( .A(arr[1930]), .B(n2646), .Y(n127) );
  AND2X1 U4238 ( .A(arr[1931]), .B(n2646), .Y(n128) );
  AND2X1 U4239 ( .A(arr[1932]), .B(n2646), .Y(n129) );
  AND2X1 U4240 ( .A(arr[1933]), .B(n2646), .Y(n130) );
  AND2X1 U4241 ( .A(arr[1934]), .B(n2646), .Y(n131) );
  AND2X1 U4242 ( .A(arr[1935]), .B(n2646), .Y(n132) );
  AND2X1 U4243 ( .A(arr[1936]), .B(n2646), .Y(n133) );
  AND2X1 U4244 ( .A(arr[1946]), .B(n2646), .Y(n134) );
  AND2X1 U4245 ( .A(arr[1952]), .B(n2645), .Y(n135) );
  AND2X1 U4246 ( .A(arr[1953]), .B(n2645), .Y(n136) );
  AND2X1 U4247 ( .A(arr[1956]), .B(n2645), .Y(n137) );
  AND2X1 U4248 ( .A(arr[1957]), .B(n2645), .Y(n138) );
  AND2X1 U4249 ( .A(arr[1958]), .B(n2645), .Y(n139) );
  AND2X1 U4250 ( .A(arr[1959]), .B(n2645), .Y(n140) );
  AND2X1 U4251 ( .A(arr[1960]), .B(n2645), .Y(n141) );
  AND2X1 U4252 ( .A(arr[1961]), .B(n2645), .Y(n142) );
  AND2X1 U4253 ( .A(arr[1962]), .B(n2645), .Y(n143) );
  AND2X1 U4254 ( .A(arr[1963]), .B(n2645), .Y(n144) );
  AND2X1 U4255 ( .A(arr[1964]), .B(n2645), .Y(n145) );
  AND2X1 U4256 ( .A(arr[1965]), .B(n2645), .Y(n146) );
  AND2X1 U4257 ( .A(arr[1966]), .B(n2645), .Y(n147) );
  AND2X1 U4258 ( .A(arr[1967]), .B(n2645), .Y(n148) );
  AND2X1 U4259 ( .A(arr[1968]), .B(n2645), .Y(n149) );
  AND2X1 U4260 ( .A(arr[1969]), .B(n2645), .Y(n150) );
  AND2X1 U4261 ( .A(arr[1979]), .B(n2645), .Y(n151) );
  AND2X1 U4262 ( .A(arr[1985]), .B(n2644), .Y(n152) );
  AND2X1 U4263 ( .A(arr[1986]), .B(n2644), .Y(n153) );
  AND2X1 U4264 ( .A(arr[1989]), .B(n2644), .Y(n154) );
  AND2X1 U4266 ( .A(arr[1990]), .B(n2644), .Y(n155) );
  AND2X1 U4267 ( .A(arr[1991]), .B(n2644), .Y(n156) );
  AND2X1 U4269 ( .A(arr[1992]), .B(n2644), .Y(n157) );
  AND2X1 U4270 ( .A(arr[1993]), .B(n2644), .Y(n158) );
  AND2X1 U4272 ( .A(arr[1994]), .B(n2644), .Y(n159) );
  AND2X1 U4273 ( .A(arr[1995]), .B(n2644), .Y(n160) );
  AND2X1 U4275 ( .A(arr[1996]), .B(n2644), .Y(n161) );
  AND2X1 U4276 ( .A(arr[1997]), .B(n2644), .Y(n162) );
  AND2X1 U4278 ( .A(arr[1998]), .B(n2644), .Y(n163) );
  AND2X1 U4279 ( .A(arr[1999]), .B(n2644), .Y(n164) );
  AND2X1 U4281 ( .A(arr[2000]), .B(n2644), .Y(n165) );
  AND2X1 U4282 ( .A(arr[2001]), .B(n2644), .Y(n166) );
  AND2X1 U4284 ( .A(arr[2002]), .B(n2644), .Y(n167) );
  AND2X1 U4285 ( .A(arr[2012]), .B(n2644), .Y(n168) );
  AND2X1 U4287 ( .A(arr[2018]), .B(n2643), .Y(n169) );
  AND2X1 U4288 ( .A(arr[2019]), .B(n2643), .Y(n170) );
  AND2X1 U4290 ( .A(arr[2022]), .B(n2643), .Y(n171) );
  AND2X1 U4291 ( .A(arr[2023]), .B(n2643), .Y(n172) );
  AND2X1 U4293 ( .A(arr[2024]), .B(n2643), .Y(n173) );
  AND2X1 U4294 ( .A(arr[2025]), .B(n2643), .Y(n174) );
  AND2X1 U4296 ( .A(arr[2026]), .B(n2643), .Y(n175) );
  AND2X1 U4297 ( .A(arr[2027]), .B(n2643), .Y(n176) );
  AND2X1 U4299 ( .A(arr[2028]), .B(n2643), .Y(n177) );
  AND2X1 U4300 ( .A(arr[2029]), .B(n2643), .Y(n178) );
  AND2X1 U4302 ( .A(arr[2030]), .B(n2643), .Y(n179) );
  AND2X1 U4303 ( .A(arr[2031]), .B(n2643), .Y(n180) );
  AND2X1 U4305 ( .A(arr[2032]), .B(n2643), .Y(n181) );
  AND2X1 U4306 ( .A(arr[2033]), .B(n2643), .Y(n182) );
  AND2X1 U4308 ( .A(arr[2034]), .B(n2643), .Y(n183) );
  AND2X1 U4309 ( .A(arr[2035]), .B(n2643), .Y(n184) );
  AND2X1 U4311 ( .A(arr[2045]), .B(n2643), .Y(n185) );
  AND2X1 U4312 ( .A(arr[2051]), .B(n2642), .Y(n186) );
  AND2X1 U4314 ( .A(arr[2052]), .B(n2642), .Y(n187) );
  AND2X1 U4315 ( .A(arr[2055]), .B(n2642), .Y(n188) );
  AND2X1 U4317 ( .A(arr[2056]), .B(n2642), .Y(n189) );
  AND2X1 U4318 ( .A(arr[2057]), .B(n2642), .Y(n190) );
  AND2X1 U4320 ( .A(arr[2058]), .B(n2642), .Y(n191) );
  AND2X1 U4321 ( .A(arr[2059]), .B(n2642), .Y(n192) );
  AND2X1 U4323 ( .A(arr[2060]), .B(n2642), .Y(n193) );
  AND2X1 U4324 ( .A(arr[2061]), .B(n2642), .Y(n194) );
  AND2X1 U4326 ( .A(arr[2062]), .B(n2642), .Y(n195) );
  AND2X1 U4327 ( .A(arr[2063]), .B(n2642), .Y(n196) );
  AND2X1 U4329 ( .A(arr[2064]), .B(n2642), .Y(n197) );
  AND2X1 U4330 ( .A(arr[2065]), .B(n2642), .Y(n198) );
  AND2X1 U4332 ( .A(arr[2066]), .B(n2642), .Y(n199) );
  AND2X1 U4333 ( .A(arr[2067]), .B(n2642), .Y(n200) );
  AND2X1 U4335 ( .A(arr[2068]), .B(n2642), .Y(n201) );
  AND2X1 U4336 ( .A(arr[2078]), .B(n2642), .Y(n202) );
  AND2X1 U4338 ( .A(arr[2084]), .B(n2641), .Y(n203) );
  AND2X1 U4339 ( .A(arr[2085]), .B(n2641), .Y(n204) );
  AND2X1 U4341 ( .A(arr[2088]), .B(n2641), .Y(n205) );
  AND2X1 U4342 ( .A(arr[2089]), .B(n2641), .Y(n206) );
  AND2X1 U4344 ( .A(arr[2090]), .B(n2641), .Y(n207) );
  AND2X1 U4345 ( .A(arr[2091]), .B(n2641), .Y(n208) );
  AND2X1 U4347 ( .A(arr[2092]), .B(n2641), .Y(n209) );
  AND2X1 U4348 ( .A(arr[2093]), .B(n2641), .Y(n210) );
  AND2X1 U4350 ( .A(arr[2094]), .B(n2641), .Y(n211) );
  AND2X1 U4351 ( .A(arr[2095]), .B(n2641), .Y(n212) );
  AND2X1 U4353 ( .A(arr[2096]), .B(n2641), .Y(n213) );
  AND2X1 U4354 ( .A(arr[2097]), .B(n2641), .Y(n214) );
  AND2X1 U4356 ( .A(arr[2098]), .B(n2641), .Y(n215) );
  AND2X1 U4357 ( .A(arr[2099]), .B(n2641), .Y(n216) );
  AND2X1 U4359 ( .A(arr[2100]), .B(n2641), .Y(n217) );
  AND2X1 U4360 ( .A(arr[2101]), .B(n2641), .Y(n218) );
  AND2X1 U4361 ( .A(arr[2111]), .B(n2641), .Y(n219) );
  AND2X1 U4365 ( .A(arr[1848]), .B(n2648), .Y(n220) );
  AND2X1 U4385 ( .A(arr[1849]), .B(n2648), .Y(n221) );
  AND2X1 U4387 ( .A(arr[1850]), .B(n2648), .Y(n222) );
  AND2X1 U4391 ( .A(arr[1851]), .B(n2648), .Y(n223) );
  AND2X1 U4431 ( .A(arr[1852]), .B(n2648), .Y(n224) );
  AND2X1 U4432 ( .A(arr[1855]), .B(n2648), .Y(n225) );
  AND2X1 U4433 ( .A(arr[1856]), .B(n2648), .Y(n226) );
  AND2X1 U4434 ( .A(arr[1871]), .B(n2648), .Y(n227) );
  AND2X1 U4435 ( .A(arr[1872]), .B(n2648), .Y(n228) );
  AND2X1 U4436 ( .A(arr[1873]), .B(n2648), .Y(n229) );
  AND2X1 U4437 ( .A(arr[1874]), .B(n2648), .Y(n230) );
  AND2X1 U4438 ( .A(arr[1875]), .B(n2648), .Y(n231) );
  AND2X1 U4439 ( .A(arr[1876]), .B(n2648), .Y(n232) );
  AND2X1 U4440 ( .A(arr[1877]), .B(n2648), .Y(n233) );
  AND2X1 U4441 ( .A(arr[1878]), .B(n2648), .Y(n234) );
  AND2X1 U4442 ( .A(arr[1879]), .B(n2648), .Y(n235) );
  AND2X1 U4443 ( .A(arr[1881]), .B(n2647), .Y(n236) );
  AND2X1 U4444 ( .A(arr[1882]), .B(n2647), .Y(n237) );
  AND2X1 U4445 ( .A(arr[1883]), .B(n2647), .Y(n238) );
  AND2X1 U4446 ( .A(arr[1884]), .B(n2647), .Y(n239) );
  AND2X1 U4447 ( .A(arr[1885]), .B(n2647), .Y(n240) );
  AND2X1 U4448 ( .A(arr[1888]), .B(n2647), .Y(n241) );
  AND2X1 U4449 ( .A(arr[1889]), .B(n2647), .Y(n242) );
  AND2X1 U4450 ( .A(arr[1904]), .B(n2647), .Y(n243) );
  AND2X1 U4451 ( .A(arr[1905]), .B(n2647), .Y(n244) );
  AND2X1 U4452 ( .A(arr[1906]), .B(n2647), .Y(n245) );
  AND2X1 U4453 ( .A(arr[1907]), .B(n2647), .Y(n246) );
  AND2X1 U4454 ( .A(arr[1908]), .B(n2647), .Y(n247) );
  AND2X1 U4455 ( .A(arr[1909]), .B(n2647), .Y(n248) );
  AND2X1 U4456 ( .A(arr[1910]), .B(n2647), .Y(n249) );
  AND2X1 U4457 ( .A(arr[1911]), .B(n2647), .Y(n250) );
  AND2X1 U4458 ( .A(arr[1912]), .B(n2647), .Y(n251) );
  AND2X1 U4459 ( .A(arr[1914]), .B(n2646), .Y(n252) );
  AND2X1 U4460 ( .A(arr[1915]), .B(n2646), .Y(n253) );
  AND2X1 U4461 ( .A(arr[1916]), .B(n2646), .Y(n254) );
  AND2X1 U4462 ( .A(arr[1917]), .B(n2646), .Y(n255) );
  AND2X1 U4463 ( .A(arr[1918]), .B(n2646), .Y(n256) );
  AND2X1 U4464 ( .A(arr[1921]), .B(n2646), .Y(n257) );
  AND2X1 U4465 ( .A(arr[1922]), .B(n2646), .Y(n258) );
  AND2X1 U4466 ( .A(arr[1937]), .B(n2646), .Y(n259) );
  AND2X1 U4467 ( .A(arr[1938]), .B(n2646), .Y(n260) );
  AND2X1 U4468 ( .A(arr[1939]), .B(n2646), .Y(n261) );
  AND2X1 U4469 ( .A(arr[1940]), .B(n2646), .Y(n262) );
  AND2X1 U4470 ( .A(arr[1941]), .B(n2646), .Y(n263) );
  AND2X1 U4471 ( .A(arr[1942]), .B(n2646), .Y(n264) );
  AND2X1 U4472 ( .A(arr[1943]), .B(n2646), .Y(n265) );
  AND2X1 U4473 ( .A(arr[1944]), .B(n2646), .Y(n266) );
  AND2X1 U4474 ( .A(arr[1945]), .B(n2646), .Y(n267) );
  AND2X1 U4475 ( .A(arr[1947]), .B(n2645), .Y(n268) );
  AND2X1 U4476 ( .A(arr[1948]), .B(n2645), .Y(n269) );
  AND2X1 U4477 ( .A(arr[1949]), .B(n2645), .Y(n270) );
  AND2X1 U4478 ( .A(arr[1950]), .B(n2645), .Y(n271) );
  AND2X1 U4479 ( .A(arr[1951]), .B(n2645), .Y(n272) );
  AND2X1 U4480 ( .A(arr[1954]), .B(n2645), .Y(n273) );
  AND2X1 U4481 ( .A(arr[1955]), .B(n2645), .Y(n274) );
  AND2X1 U4482 ( .A(arr[1970]), .B(n2645), .Y(n275) );
  AND2X1 U4483 ( .A(arr[1971]), .B(n2645), .Y(n276) );
  AND2X1 U4484 ( .A(arr[1972]), .B(n2645), .Y(n277) );
  AND2X1 U4485 ( .A(arr[1973]), .B(n2645), .Y(n278) );
  AND2X1 U4486 ( .A(arr[1974]), .B(n2645), .Y(n279) );
  AND2X1 U4487 ( .A(arr[1975]), .B(n2645), .Y(n280) );
  AND2X1 U4488 ( .A(arr[1976]), .B(n2645), .Y(n281) );
  AND2X1 U4489 ( .A(arr[1977]), .B(n2645), .Y(n282) );
  AND2X1 U4490 ( .A(arr[1978]), .B(n2645), .Y(n283) );
  AND2X1 U4491 ( .A(arr[1980]), .B(n2644), .Y(n284) );
  AND2X1 U4492 ( .A(arr[1981]), .B(n2644), .Y(n285) );
  AND2X1 U4493 ( .A(arr[1982]), .B(n2644), .Y(n286) );
  AND2X1 U4494 ( .A(arr[1983]), .B(n2644), .Y(n287) );
  AND2X1 U4495 ( .A(arr[1984]), .B(n2644), .Y(n288) );
  AND2X1 U4496 ( .A(arr[1987]), .B(n2644), .Y(n289) );
  AND2X1 U4497 ( .A(arr[1988]), .B(n2644), .Y(n290) );
  AND2X1 U4498 ( .A(arr[2003]), .B(n2644), .Y(n291) );
  AND2X1 U4499 ( .A(arr[2004]), .B(n2644), .Y(n292) );
  AND2X1 U4500 ( .A(arr[2005]), .B(n2644), .Y(n293) );
  AND2X1 U4501 ( .A(arr[2006]), .B(n2644), .Y(n294) );
  AND2X1 U4502 ( .A(arr[2007]), .B(n2644), .Y(n295) );
  AND2X1 U4503 ( .A(arr[2008]), .B(n2644), .Y(n296) );
  AND2X1 U4504 ( .A(arr[2009]), .B(n2644), .Y(n297) );
  AND2X1 U4505 ( .A(arr[2010]), .B(n2644), .Y(n298) );
  AND2X1 U4506 ( .A(arr[2011]), .B(n2644), .Y(n299) );
  AND2X1 U4507 ( .A(arr[2013]), .B(n2643), .Y(n300) );
  AND2X1 U4508 ( .A(arr[2014]), .B(n2643), .Y(n301) );
  AND2X1 U4509 ( .A(arr[2015]), .B(n2643), .Y(n302) );
  AND2X1 U4510 ( .A(arr[2016]), .B(n2643), .Y(n303) );
  AND2X1 U4511 ( .A(arr[2017]), .B(n2643), .Y(n304) );
  AND2X1 U4512 ( .A(arr[2020]), .B(n2643), .Y(n305) );
  AND2X1 U4513 ( .A(arr[2021]), .B(n2643), .Y(n306) );
  AND2X1 U4514 ( .A(arr[2036]), .B(n2643), .Y(n307) );
  AND2X1 U4515 ( .A(arr[2037]), .B(n2643), .Y(n308) );
  AND2X1 U4516 ( .A(arr[2038]), .B(n2643), .Y(n309) );
  AND2X1 U4517 ( .A(arr[2039]), .B(n2643), .Y(n310) );
  AND2X1 U4518 ( .A(arr[2040]), .B(n2643), .Y(n311) );
  AND2X1 U4519 ( .A(arr[2041]), .B(n2643), .Y(n312) );
  AND2X1 U4520 ( .A(arr[2042]), .B(n2643), .Y(n313) );
  AND2X1 U4521 ( .A(arr[2043]), .B(n2643), .Y(n314) );
  AND2X1 U4522 ( .A(arr[2044]), .B(n2643), .Y(n315) );
  AND2X1 U4523 ( .A(arr[2046]), .B(n2642), .Y(n316) );
  AND2X1 U4524 ( .A(arr[2047]), .B(n2642), .Y(n317) );
  AND2X1 U4525 ( .A(arr[2048]), .B(n2642), .Y(n318) );
  AND2X1 U4526 ( .A(arr[2049]), .B(n2642), .Y(n319) );
  AND2X1 U4527 ( .A(arr[2050]), .B(n2642), .Y(n320) );
  AND2X1 U4528 ( .A(arr[2053]), .B(n2642), .Y(n321) );
  AND2X1 U4529 ( .A(arr[2054]), .B(n2642), .Y(n322) );
  AND2X1 U4530 ( .A(arr[2069]), .B(n2642), .Y(n323) );
  AND2X1 U4531 ( .A(arr[2070]), .B(n2642), .Y(n324) );
  AND2X1 U4532 ( .A(arr[2071]), .B(n2642), .Y(n325) );
  AND2X1 U4533 ( .A(arr[2072]), .B(n2642), .Y(n326) );
  AND2X1 U4534 ( .A(arr[2073]), .B(n2642), .Y(n327) );
  AND2X1 U4535 ( .A(arr[2074]), .B(n2642), .Y(n328) );
  AND2X1 U4536 ( .A(arr[2075]), .B(n2642), .Y(n329) );
  AND2X1 U4537 ( .A(arr[2076]), .B(n2642), .Y(n330) );
  AND2X1 U4538 ( .A(arr[2077]), .B(n2642), .Y(n331) );
  AND2X1 U4539 ( .A(arr[2079]), .B(n2641), .Y(n332) );
  AND2X1 U4540 ( .A(arr[2080]), .B(n2641), .Y(n333) );
  AND2X1 U4541 ( .A(arr[2081]), .B(n2641), .Y(n334) );
  AND2X1 U4542 ( .A(arr[2082]), .B(n2641), .Y(n335) );
  AND2X1 U4543 ( .A(arr[2083]), .B(n2641), .Y(n336) );
  AND2X1 U4544 ( .A(arr[2086]), .B(n2641), .Y(n337) );
  AND2X1 U4545 ( .A(arr[2087]), .B(n2641), .Y(n338) );
  AND2X1 U4546 ( .A(arr[2102]), .B(n2641), .Y(n339) );
  AND2X1 U4547 ( .A(arr[2103]), .B(n2641), .Y(n340) );
  AND2X1 U4548 ( .A(arr[2104]), .B(n2641), .Y(n341) );
  AND2X1 U4549 ( .A(arr[2105]), .B(n2641), .Y(n342) );
  AND2X1 U4550 ( .A(arr[2106]), .B(n2641), .Y(n343) );
  AND2X1 U4551 ( .A(arr[2107]), .B(n2641), .Y(n344) );
  AND2X1 U4552 ( .A(arr[2108]), .B(n2641), .Y(n345) );
  AND2X1 U4553 ( .A(arr[2109]), .B(n2641), .Y(n346) );
  AND2X1 U4554 ( .A(arr[2110]), .B(n2641), .Y(n347) );
  BUFX2 U4555 ( .A(n2616), .Y(n2594) );
  BUFX2 U4556 ( .A(n15), .Y(n2616) );
  BUFX2 U4557 ( .A(n17), .Y(n2636) );
  BUFX2 U4558 ( .A(n17), .Y(n2637) );
  BUFX2 U4559 ( .A(n17), .Y(n2638) );
  BUFX2 U4560 ( .A(n17), .Y(n2639) );
  BUFX2 U4561 ( .A(n17), .Y(n2640) );
  BUFX2 U4562 ( .A(n17), .Y(n2635) );
  BUFX2 U4563 ( .A(n15), .Y(n2617) );
  BUFX2 U4564 ( .A(n15), .Y(n2618) );
  BUFX2 U4565 ( .A(n15), .Y(n2619) );
  BUFX2 U4566 ( .A(n15), .Y(n2620) );
  BUFX2 U4567 ( .A(n15), .Y(n2621) );
  BUFX2 U4568 ( .A(n15), .Y(n2622) );
  BUFX2 U4569 ( .A(n15), .Y(n2623) );
  MUX2X1 U4570 ( .B(n349), .A(n350), .S(n2535), .Y(n348) );
  MUX2X1 U4571 ( .B(n352), .A(n353), .S(n2535), .Y(n351) );
  MUX2X1 U4572 ( .B(n355), .A(n356), .S(n2535), .Y(n354) );
  MUX2X1 U4573 ( .B(n358), .A(n359), .S(n2535), .Y(n357) );
  MUX2X1 U4574 ( .B(n361), .A(n362), .S(n2624), .Y(n360) );
  MUX2X1 U4575 ( .B(n364), .A(n365), .S(n2535), .Y(n363) );
  MUX2X1 U4576 ( .B(n367), .A(n368), .S(n2535), .Y(n366) );
  MUX2X1 U4577 ( .B(n370), .A(n371), .S(n2535), .Y(n369) );
  MUX2X1 U4578 ( .B(n373), .A(n374), .S(n2535), .Y(n372) );
  MUX2X1 U4579 ( .B(n376), .A(n377), .S(n2624), .Y(n375) );
  MUX2X1 U4580 ( .B(n379), .A(n380), .S(n2535), .Y(n378) );
  MUX2X1 U4581 ( .B(n382), .A(n383), .S(n2535), .Y(n381) );
  MUX2X1 U4582 ( .B(n385), .A(n386), .S(n2535), .Y(n384) );
  MUX2X1 U4583 ( .B(n388), .A(n389), .S(n2535), .Y(n387) );
  MUX2X1 U4584 ( .B(n391), .A(n392), .S(n2624), .Y(n390) );
  MUX2X1 U4585 ( .B(n394), .A(n395), .S(n2536), .Y(n393) );
  MUX2X1 U4586 ( .B(n397), .A(n398), .S(n2536), .Y(n396) );
  MUX2X1 U4587 ( .B(n400), .A(n401), .S(n2536), .Y(n399) );
  MUX2X1 U4588 ( .B(n403), .A(n404), .S(n2536), .Y(n402) );
  MUX2X1 U4589 ( .B(n406), .A(n407), .S(n2624), .Y(n405) );
  MUX2X1 U4590 ( .B(n408), .A(n409), .S(n18), .Y(data_out[0]) );
  MUX2X1 U4591 ( .B(n411), .A(n412), .S(n2536), .Y(n410) );
  MUX2X1 U4592 ( .B(n414), .A(n415), .S(n2536), .Y(n413) );
  MUX2X1 U4593 ( .B(n417), .A(n418), .S(n2536), .Y(n416) );
  MUX2X1 U4594 ( .B(n420), .A(n421), .S(n2536), .Y(n419) );
  MUX2X1 U4595 ( .B(n423), .A(n424), .S(n2624), .Y(n422) );
  MUX2X1 U4596 ( .B(n426), .A(n427), .S(n2536), .Y(n425) );
  MUX2X1 U4597 ( .B(n429), .A(n430), .S(n2536), .Y(n428) );
  MUX2X1 U4598 ( .B(n432), .A(n433), .S(n2536), .Y(n431) );
  MUX2X1 U4599 ( .B(n435), .A(n436), .S(n2536), .Y(n434) );
  MUX2X1 U4600 ( .B(n438), .A(n439), .S(n2624), .Y(n437) );
  MUX2X1 U4601 ( .B(n441), .A(n442), .S(n2537), .Y(n440) );
  MUX2X1 U4602 ( .B(n444), .A(n445), .S(n2537), .Y(n443) );
  MUX2X1 U4603 ( .B(n447), .A(n448), .S(n2537), .Y(n446) );
  MUX2X1 U4604 ( .B(n450), .A(n451), .S(n2537), .Y(n449) );
  MUX2X1 U4605 ( .B(n453), .A(n454), .S(n2624), .Y(n452) );
  MUX2X1 U4606 ( .B(n456), .A(n457), .S(n2537), .Y(n455) );
  MUX2X1 U4607 ( .B(n459), .A(n460), .S(n2537), .Y(n458) );
  MUX2X1 U4608 ( .B(n462), .A(n463), .S(n2537), .Y(n461) );
  MUX2X1 U4609 ( .B(n465), .A(n466), .S(n2537), .Y(n464) );
  MUX2X1 U4610 ( .B(n468), .A(n469), .S(n2624), .Y(n467) );
  MUX2X1 U4611 ( .B(n470), .A(n471), .S(n18), .Y(data_out[1]) );
  MUX2X1 U4612 ( .B(n473), .A(n474), .S(n2537), .Y(n472) );
  MUX2X1 U4613 ( .B(n476), .A(n477), .S(n2537), .Y(n475) );
  MUX2X1 U4614 ( .B(n479), .A(n480), .S(n2537), .Y(n478) );
  MUX2X1 U4615 ( .B(n482), .A(n483), .S(n2537), .Y(n481) );
  MUX2X1 U4616 ( .B(n485), .A(n486), .S(n2624), .Y(n484) );
  MUX2X1 U4617 ( .B(n488), .A(n489), .S(n2538), .Y(n487) );
  MUX2X1 U4618 ( .B(n491), .A(n492), .S(n2538), .Y(n490) );
  MUX2X1 U4619 ( .B(n494), .A(n495), .S(n2538), .Y(n493) );
  MUX2X1 U4620 ( .B(n497), .A(n498), .S(n2538), .Y(n496) );
  MUX2X1 U4621 ( .B(n500), .A(n501), .S(n2624), .Y(n499) );
  MUX2X1 U4622 ( .B(n503), .A(n504), .S(n2538), .Y(n502) );
  MUX2X1 U4623 ( .B(n506), .A(n507), .S(n2538), .Y(n505) );
  MUX2X1 U4624 ( .B(n509), .A(n510), .S(n2538), .Y(n508) );
  MUX2X1 U4625 ( .B(n512), .A(n513), .S(n2538), .Y(n511) );
  MUX2X1 U4626 ( .B(n515), .A(n516), .S(n2624), .Y(n514) );
  MUX2X1 U4627 ( .B(n518), .A(n519), .S(n2538), .Y(n517) );
  MUX2X1 U4628 ( .B(n521), .A(n522), .S(n2538), .Y(n520) );
  MUX2X1 U4629 ( .B(n524), .A(n525), .S(n2538), .Y(n523) );
  MUX2X1 U4630 ( .B(n527), .A(n528), .S(n2538), .Y(n526) );
  MUX2X1 U4631 ( .B(n530), .A(n531), .S(n2624), .Y(n529) );
  MUX2X1 U4632 ( .B(n532), .A(n533), .S(n18), .Y(data_out[2]) );
  MUX2X1 U4633 ( .B(n535), .A(n536), .S(n2539), .Y(n534) );
  MUX2X1 U4634 ( .B(n538), .A(n539), .S(n2539), .Y(n537) );
  MUX2X1 U4635 ( .B(n541), .A(n542), .S(n2539), .Y(n540) );
  MUX2X1 U4636 ( .B(n544), .A(n545), .S(n2539), .Y(n543) );
  MUX2X1 U4637 ( .B(n547), .A(n548), .S(n2625), .Y(n546) );
  MUX2X1 U4638 ( .B(n550), .A(n551), .S(n2539), .Y(n549) );
  MUX2X1 U4639 ( .B(n553), .A(n554), .S(n2539), .Y(n552) );
  MUX2X1 U4640 ( .B(n556), .A(n557), .S(n2539), .Y(n555) );
  MUX2X1 U4641 ( .B(n559), .A(n560), .S(n2539), .Y(n558) );
  MUX2X1 U4642 ( .B(n562), .A(n563), .S(n2625), .Y(n561) );
  MUX2X1 U4643 ( .B(n565), .A(n566), .S(n2539), .Y(n564) );
  MUX2X1 U4644 ( .B(n568), .A(n569), .S(n2539), .Y(n567) );
  MUX2X1 U4645 ( .B(n571), .A(n572), .S(n2539), .Y(n570) );
  MUX2X1 U4646 ( .B(n574), .A(n575), .S(n2539), .Y(n573) );
  MUX2X1 U4647 ( .B(n577), .A(n578), .S(n2625), .Y(n576) );
  MUX2X1 U4648 ( .B(n580), .A(n581), .S(n2540), .Y(n579) );
  MUX2X1 U4649 ( .B(n583), .A(n584), .S(n2540), .Y(n582) );
  MUX2X1 U4650 ( .B(n586), .A(n587), .S(n2540), .Y(n585) );
  MUX2X1 U4651 ( .B(n589), .A(n590), .S(n2540), .Y(n588) );
  MUX2X1 U4652 ( .B(n592), .A(n593), .S(n2625), .Y(n591) );
  MUX2X1 U4653 ( .B(n594), .A(n595), .S(n18), .Y(data_out[3]) );
  MUX2X1 U4654 ( .B(n597), .A(n598), .S(n2540), .Y(n596) );
  MUX2X1 U4655 ( .B(n600), .A(n601), .S(n2540), .Y(n599) );
  MUX2X1 U4656 ( .B(n603), .A(n604), .S(n2540), .Y(n602) );
  MUX2X1 U4657 ( .B(n606), .A(n607), .S(n2540), .Y(n605) );
  MUX2X1 U4658 ( .B(n609), .A(n610), .S(n2625), .Y(n608) );
  MUX2X1 U4659 ( .B(n612), .A(n613), .S(n2540), .Y(n611) );
  MUX2X1 U4660 ( .B(n615), .A(n616), .S(n2540), .Y(n614) );
  MUX2X1 U4661 ( .B(n618), .A(n619), .S(n2540), .Y(n617) );
  MUX2X1 U4662 ( .B(n621), .A(n622), .S(n2540), .Y(n620) );
  MUX2X1 U4663 ( .B(n624), .A(n625), .S(n2625), .Y(n623) );
  MUX2X1 U4664 ( .B(n627), .A(n628), .S(n2541), .Y(n626) );
  MUX2X1 U4665 ( .B(n630), .A(n631), .S(n2541), .Y(n629) );
  MUX2X1 U4666 ( .B(n633), .A(n634), .S(n2541), .Y(n632) );
  MUX2X1 U4667 ( .B(n636), .A(n637), .S(n2541), .Y(n635) );
  MUX2X1 U4668 ( .B(n639), .A(n640), .S(n2625), .Y(n638) );
  MUX2X1 U4669 ( .B(n642), .A(n643), .S(n2541), .Y(n641) );
  MUX2X1 U4670 ( .B(n645), .A(n646), .S(n2541), .Y(n644) );
  MUX2X1 U4671 ( .B(n648), .A(n649), .S(n2541), .Y(n647) );
  MUX2X1 U4672 ( .B(n651), .A(n652), .S(n2541), .Y(n650) );
  MUX2X1 U4673 ( .B(n654), .A(n655), .S(n2625), .Y(n653) );
  MUX2X1 U4674 ( .B(n656), .A(n657), .S(n18), .Y(data_out[4]) );
  MUX2X1 U4675 ( .B(n659), .A(n660), .S(n2541), .Y(n658) );
  MUX2X1 U4676 ( .B(n662), .A(n663), .S(n2541), .Y(n661) );
  MUX2X1 U4677 ( .B(n665), .A(n666), .S(n2541), .Y(n664) );
  MUX2X1 U4678 ( .B(n668), .A(n669), .S(n2541), .Y(n667) );
  MUX2X1 U4679 ( .B(n671), .A(n672), .S(n2625), .Y(n670) );
  MUX2X1 U4680 ( .B(n674), .A(n675), .S(n2542), .Y(n673) );
  MUX2X1 U4681 ( .B(n677), .A(n678), .S(n2542), .Y(n676) );
  MUX2X1 U4682 ( .B(n680), .A(n681), .S(n2542), .Y(n679) );
  MUX2X1 U4683 ( .B(n683), .A(n684), .S(n2542), .Y(n682) );
  MUX2X1 U4684 ( .B(n686), .A(n687), .S(n2625), .Y(n685) );
  MUX2X1 U4685 ( .B(n689), .A(n690), .S(n2542), .Y(n688) );
  MUX2X1 U4686 ( .B(n692), .A(n693), .S(n2542), .Y(n691) );
  MUX2X1 U4687 ( .B(n695), .A(n696), .S(n2542), .Y(n694) );
  MUX2X1 U4688 ( .B(n698), .A(n699), .S(n2542), .Y(n697) );
  MUX2X1 U4689 ( .B(n701), .A(n702), .S(n2625), .Y(n700) );
  MUX2X1 U4690 ( .B(n704), .A(n705), .S(n2542), .Y(n703) );
  MUX2X1 U4691 ( .B(n707), .A(n708), .S(n2542), .Y(n706) );
  MUX2X1 U4692 ( .B(n710), .A(n711), .S(n2542), .Y(n709) );
  MUX2X1 U4693 ( .B(n713), .A(n714), .S(n2542), .Y(n712) );
  MUX2X1 U4694 ( .B(n716), .A(n717), .S(n2625), .Y(n715) );
  MUX2X1 U4695 ( .B(n718), .A(n719), .S(n18), .Y(data_out[5]) );
  MUX2X1 U4696 ( .B(n721), .A(n722), .S(n2543), .Y(n720) );
  MUX2X1 U4697 ( .B(n724), .A(n725), .S(n2543), .Y(n723) );
  MUX2X1 U4698 ( .B(n727), .A(n728), .S(n2543), .Y(n726) );
  MUX2X1 U4699 ( .B(n730), .A(n731), .S(n2543), .Y(n729) );
  MUX2X1 U4700 ( .B(n733), .A(n734), .S(n2626), .Y(n732) );
  MUX2X1 U4701 ( .B(n736), .A(n737), .S(n2543), .Y(n735) );
  MUX2X1 U4702 ( .B(n739), .A(n740), .S(n2543), .Y(n738) );
  MUX2X1 U4703 ( .B(n742), .A(n743), .S(n2543), .Y(n741) );
  MUX2X1 U4704 ( .B(n745), .A(n746), .S(n2543), .Y(n744) );
  MUX2X1 U4705 ( .B(n748), .A(n749), .S(n2626), .Y(n747) );
  MUX2X1 U4706 ( .B(n751), .A(n752), .S(n2543), .Y(n750) );
  MUX2X1 U4707 ( .B(n754), .A(n755), .S(n2543), .Y(n753) );
  MUX2X1 U4708 ( .B(n757), .A(n758), .S(n2543), .Y(n756) );
  MUX2X1 U4709 ( .B(n760), .A(n761), .S(n2543), .Y(n759) );
  MUX2X1 U4710 ( .B(n763), .A(n764), .S(n2626), .Y(n762) );
  MUX2X1 U4711 ( .B(n766), .A(n767), .S(n2544), .Y(n765) );
  MUX2X1 U4712 ( .B(n769), .A(n770), .S(n2544), .Y(n768) );
  MUX2X1 U4713 ( .B(n772), .A(n773), .S(n2544), .Y(n771) );
  MUX2X1 U4714 ( .B(n775), .A(n776), .S(n2544), .Y(n774) );
  MUX2X1 U4715 ( .B(n778), .A(n779), .S(n2626), .Y(n777) );
  MUX2X1 U4716 ( .B(n780), .A(n781), .S(n18), .Y(data_out[6]) );
  MUX2X1 U4717 ( .B(n783), .A(n784), .S(n2544), .Y(n782) );
  MUX2X1 U4718 ( .B(n786), .A(n787), .S(n2544), .Y(n785) );
  MUX2X1 U4719 ( .B(n789), .A(n790), .S(n2544), .Y(n788) );
  MUX2X1 U4720 ( .B(n792), .A(n793), .S(n2544), .Y(n791) );
  MUX2X1 U4721 ( .B(n795), .A(n796), .S(n2626), .Y(n794) );
  MUX2X1 U4722 ( .B(n798), .A(n799), .S(n2544), .Y(n797) );
  MUX2X1 U4723 ( .B(n801), .A(n802), .S(n2544), .Y(n800) );
  MUX2X1 U4724 ( .B(n804), .A(n805), .S(n2544), .Y(n803) );
  MUX2X1 U4725 ( .B(n807), .A(n808), .S(n2544), .Y(n806) );
  MUX2X1 U4726 ( .B(n810), .A(n811), .S(n2626), .Y(n809) );
  MUX2X1 U4727 ( .B(n813), .A(n814), .S(n2545), .Y(n812) );
  MUX2X1 U4728 ( .B(n816), .A(n817), .S(n2545), .Y(n815) );
  MUX2X1 U4729 ( .B(n819), .A(n820), .S(n2545), .Y(n818) );
  MUX2X1 U4730 ( .B(n822), .A(n823), .S(n2545), .Y(n821) );
  MUX2X1 U4731 ( .B(n825), .A(n826), .S(n2626), .Y(n824) );
  MUX2X1 U4732 ( .B(n828), .A(n829), .S(n2545), .Y(n827) );
  MUX2X1 U4733 ( .B(n831), .A(n832), .S(n2545), .Y(n830) );
  MUX2X1 U4734 ( .B(n834), .A(n835), .S(n2545), .Y(n833) );
  MUX2X1 U4735 ( .B(n837), .A(n838), .S(n2545), .Y(n836) );
  MUX2X1 U4736 ( .B(n840), .A(n841), .S(n2626), .Y(n839) );
  MUX2X1 U4737 ( .B(n842), .A(n843), .S(n18), .Y(data_out[7]) );
  MUX2X1 U4738 ( .B(n845), .A(n846), .S(n2545), .Y(n844) );
  MUX2X1 U4739 ( .B(n848), .A(n849), .S(n2545), .Y(n847) );
  MUX2X1 U4740 ( .B(n851), .A(n852), .S(n2545), .Y(n850) );
  MUX2X1 U4741 ( .B(n854), .A(n855), .S(n2545), .Y(n853) );
  MUX2X1 U4742 ( .B(n857), .A(n858), .S(n2626), .Y(n856) );
  MUX2X1 U4743 ( .B(n860), .A(n861), .S(n2546), .Y(n859) );
  MUX2X1 U4744 ( .B(n863), .A(n864), .S(n2546), .Y(n862) );
  MUX2X1 U4745 ( .B(n866), .A(n867), .S(n2546), .Y(n865) );
  MUX2X1 U4746 ( .B(n869), .A(n870), .S(n2546), .Y(n868) );
  MUX2X1 U4747 ( .B(n872), .A(n873), .S(n2626), .Y(n871) );
  MUX2X1 U4748 ( .B(n875), .A(n876), .S(n2546), .Y(n874) );
  MUX2X1 U4749 ( .B(n878), .A(n879), .S(n2546), .Y(n877) );
  MUX2X1 U4750 ( .B(n881), .A(n882), .S(n2546), .Y(n880) );
  MUX2X1 U4751 ( .B(n884), .A(n885), .S(n2546), .Y(n883) );
  MUX2X1 U4752 ( .B(n887), .A(n888), .S(n2626), .Y(n886) );
  MUX2X1 U4753 ( .B(n890), .A(n891), .S(n2546), .Y(n889) );
  MUX2X1 U4754 ( .B(n893), .A(n894), .S(n2546), .Y(n892) );
  MUX2X1 U4755 ( .B(n896), .A(n897), .S(n2546), .Y(n895) );
  MUX2X1 U4756 ( .B(n899), .A(n900), .S(n2546), .Y(n898) );
  MUX2X1 U4757 ( .B(n902), .A(n903), .S(n2626), .Y(n901) );
  MUX2X1 U4758 ( .B(n904), .A(n905), .S(n18), .Y(data_out[8]) );
  MUX2X1 U4759 ( .B(n907), .A(n908), .S(n2547), .Y(n906) );
  MUX2X1 U4760 ( .B(n910), .A(n911), .S(n2547), .Y(n909) );
  MUX2X1 U4761 ( .B(n913), .A(n914), .S(n2547), .Y(n912) );
  MUX2X1 U4762 ( .B(n916), .A(n917), .S(n2547), .Y(n915) );
  MUX2X1 U4763 ( .B(n919), .A(n920), .S(n2627), .Y(n918) );
  MUX2X1 U4764 ( .B(n922), .A(n923), .S(n2547), .Y(n921) );
  MUX2X1 U4765 ( .B(n925), .A(n926), .S(n2547), .Y(n924) );
  MUX2X1 U4766 ( .B(n928), .A(n929), .S(n2547), .Y(n927) );
  MUX2X1 U4767 ( .B(n931), .A(n932), .S(n2547), .Y(n930) );
  MUX2X1 U4768 ( .B(n934), .A(n935), .S(n2627), .Y(n933) );
  MUX2X1 U4769 ( .B(n937), .A(n938), .S(n2547), .Y(n936) );
  MUX2X1 U4770 ( .B(n940), .A(n941), .S(n2547), .Y(n939) );
  MUX2X1 U4771 ( .B(n943), .A(n944), .S(n2547), .Y(n942) );
  MUX2X1 U4772 ( .B(n946), .A(n947), .S(n2547), .Y(n945) );
  MUX2X1 U4773 ( .B(n949), .A(n950), .S(n2627), .Y(n948) );
  MUX2X1 U4774 ( .B(n952), .A(n953), .S(n2548), .Y(n951) );
  MUX2X1 U4775 ( .B(n955), .A(n956), .S(n2548), .Y(n954) );
  MUX2X1 U4776 ( .B(n958), .A(n959), .S(n2548), .Y(n957) );
  MUX2X1 U4777 ( .B(n961), .A(n962), .S(n2548), .Y(n960) );
  MUX2X1 U4778 ( .B(n964), .A(n965), .S(n2627), .Y(n963) );
  MUX2X1 U4779 ( .B(n966), .A(n967), .S(n18), .Y(data_out[9]) );
  MUX2X1 U4780 ( .B(n969), .A(n970), .S(n2548), .Y(n968) );
  MUX2X1 U4781 ( .B(n972), .A(n973), .S(n2548), .Y(n971) );
  MUX2X1 U4782 ( .B(n975), .A(n976), .S(n2548), .Y(n974) );
  MUX2X1 U4783 ( .B(n978), .A(n979), .S(n2548), .Y(n977) );
  MUX2X1 U4784 ( .B(n981), .A(n982), .S(n2627), .Y(n980) );
  MUX2X1 U4785 ( .B(n984), .A(n985), .S(n2548), .Y(n983) );
  MUX2X1 U4786 ( .B(n987), .A(n988), .S(n2548), .Y(n986) );
  MUX2X1 U4787 ( .B(n990), .A(n991), .S(n2548), .Y(n989) );
  MUX2X1 U4788 ( .B(n993), .A(n994), .S(n2548), .Y(n992) );
  MUX2X1 U4789 ( .B(n996), .A(n997), .S(n2627), .Y(n995) );
  MUX2X1 U4790 ( .B(n999), .A(n1000), .S(n2549), .Y(n998) );
  MUX2X1 U4791 ( .B(n1002), .A(n1003), .S(n2549), .Y(n1001) );
  MUX2X1 U4792 ( .B(n1005), .A(n1006), .S(n2549), .Y(n1004) );
  MUX2X1 U4793 ( .B(n1008), .A(n1009), .S(n2549), .Y(n1007) );
  MUX2X1 U4794 ( .B(n1011), .A(n1012), .S(n2627), .Y(n1010) );
  MUX2X1 U4795 ( .B(n1014), .A(n1015), .S(n2549), .Y(n1013) );
  MUX2X1 U4796 ( .B(n1017), .A(n1018), .S(n2549), .Y(n1016) );
  MUX2X1 U4797 ( .B(n1020), .A(n1021), .S(n2549), .Y(n1019) );
  MUX2X1 U4798 ( .B(n1023), .A(n1024), .S(n2549), .Y(n1022) );
  MUX2X1 U4799 ( .B(n1026), .A(n1027), .S(n2627), .Y(n1025) );
  MUX2X1 U4800 ( .B(n1028), .A(n1029), .S(n18), .Y(data_out[10]) );
  MUX2X1 U4801 ( .B(n1031), .A(n1032), .S(n2549), .Y(n1030) );
  MUX2X1 U4802 ( .B(n1034), .A(n1035), .S(n2549), .Y(n1033) );
  MUX2X1 U4803 ( .B(n1037), .A(n1038), .S(n2549), .Y(n1036) );
  MUX2X1 U4804 ( .B(n1040), .A(n1041), .S(n2549), .Y(n1039) );
  MUX2X1 U4805 ( .B(n1043), .A(n1044), .S(n2627), .Y(n1042) );
  MUX2X1 U4806 ( .B(n1046), .A(n1047), .S(n2550), .Y(n1045) );
  MUX2X1 U4807 ( .B(n1049), .A(n1050), .S(n2550), .Y(n1048) );
  MUX2X1 U4808 ( .B(n1052), .A(n1053), .S(n2550), .Y(n1051) );
  MUX2X1 U4809 ( .B(n1055), .A(n1056), .S(n2550), .Y(n1054) );
  MUX2X1 U4810 ( .B(n1058), .A(n1059), .S(n2627), .Y(n1057) );
  MUX2X1 U4811 ( .B(n1061), .A(n1062), .S(n2550), .Y(n1060) );
  MUX2X1 U4812 ( .B(n1064), .A(n1065), .S(n2550), .Y(n1063) );
  MUX2X1 U4813 ( .B(n1067), .A(n1068), .S(n2550), .Y(n1066) );
  MUX2X1 U4814 ( .B(n1070), .A(n1071), .S(n2550), .Y(n1069) );
  MUX2X1 U4815 ( .B(n1073), .A(n1074), .S(n2627), .Y(n1072) );
  MUX2X1 U4816 ( .B(n1076), .A(n1077), .S(n2550), .Y(n1075) );
  MUX2X1 U4817 ( .B(n1079), .A(n1080), .S(n2550), .Y(n1078) );
  MUX2X1 U4818 ( .B(n1082), .A(n1083), .S(n2550), .Y(n1081) );
  MUX2X1 U4819 ( .B(n1085), .A(n1086), .S(n2550), .Y(n1084) );
  MUX2X1 U4820 ( .B(n1088), .A(n1089), .S(n2627), .Y(n1087) );
  MUX2X1 U4821 ( .B(n1090), .A(n1091), .S(n18), .Y(data_out[11]) );
  MUX2X1 U4822 ( .B(n1093), .A(n1094), .S(n2551), .Y(n1092) );
  MUX2X1 U4823 ( .B(n1096), .A(n1097), .S(n2551), .Y(n1095) );
  MUX2X1 U4824 ( .B(n1099), .A(n1100), .S(n2551), .Y(n1098) );
  MUX2X1 U4825 ( .B(n1102), .A(n1103), .S(n2551), .Y(n1101) );
  MUX2X1 U4826 ( .B(n1105), .A(n1106), .S(n2628), .Y(n1104) );
  MUX2X1 U4827 ( .B(n1108), .A(n1109), .S(n2551), .Y(n1107) );
  MUX2X1 U4828 ( .B(n1111), .A(n1112), .S(n2551), .Y(n1110) );
  MUX2X1 U4829 ( .B(n1114), .A(n1115), .S(n2551), .Y(n1113) );
  MUX2X1 U4830 ( .B(n1117), .A(n1118), .S(n2551), .Y(n1116) );
  MUX2X1 U4831 ( .B(n1120), .A(n1121), .S(n2628), .Y(n1119) );
  MUX2X1 U4832 ( .B(n1123), .A(n1124), .S(n2551), .Y(n1122) );
  MUX2X1 U4833 ( .B(n1126), .A(n1127), .S(n2551), .Y(n1125) );
  MUX2X1 U4834 ( .B(n1129), .A(n1130), .S(n2551), .Y(n1128) );
  MUX2X1 U4835 ( .B(n1132), .A(n1133), .S(n2551), .Y(n1131) );
  MUX2X1 U4836 ( .B(n1135), .A(n1136), .S(n2628), .Y(n1134) );
  MUX2X1 U4837 ( .B(n1138), .A(n1139), .S(n2552), .Y(n1137) );
  MUX2X1 U4838 ( .B(n1141), .A(n1142), .S(n2552), .Y(n1140) );
  MUX2X1 U4839 ( .B(n1144), .A(n1145), .S(n2552), .Y(n1143) );
  MUX2X1 U4840 ( .B(n1147), .A(n1148), .S(n2552), .Y(n1146) );
  MUX2X1 U4841 ( .B(n1150), .A(n1151), .S(n2628), .Y(n1149) );
  MUX2X1 U4842 ( .B(n1152), .A(n1153), .S(n18), .Y(data_out[12]) );
  MUX2X1 U4843 ( .B(n1155), .A(n1156), .S(n2552), .Y(n1154) );
  MUX2X1 U4844 ( .B(n1158), .A(n1159), .S(n2552), .Y(n1157) );
  MUX2X1 U4845 ( .B(n1161), .A(n1162), .S(n2552), .Y(n1160) );
  MUX2X1 U4846 ( .B(n1164), .A(n1165), .S(n2552), .Y(n1163) );
  MUX2X1 U4847 ( .B(n1167), .A(n1168), .S(n2628), .Y(n1166) );
  MUX2X1 U4848 ( .B(n1170), .A(n1171), .S(n2552), .Y(n1169) );
  MUX2X1 U4849 ( .B(n1173), .A(n1174), .S(n2552), .Y(n1172) );
  MUX2X1 U4850 ( .B(n1176), .A(n1177), .S(n2552), .Y(n1175) );
  MUX2X1 U4851 ( .B(n1179), .A(n1180), .S(n2552), .Y(n1178) );
  MUX2X1 U4852 ( .B(n1182), .A(n1183), .S(n2628), .Y(n1181) );
  MUX2X1 U4853 ( .B(n1185), .A(n1186), .S(n2553), .Y(n1184) );
  MUX2X1 U4854 ( .B(n1188), .A(n1189), .S(n2553), .Y(n1187) );
  MUX2X1 U4855 ( .B(n1191), .A(n1192), .S(n2553), .Y(n1190) );
  MUX2X1 U4856 ( .B(n1194), .A(n1195), .S(n2553), .Y(n1193) );
  MUX2X1 U4857 ( .B(n1197), .A(n1198), .S(n2628), .Y(n1196) );
  MUX2X1 U4858 ( .B(n1200), .A(n1201), .S(n2553), .Y(n1199) );
  MUX2X1 U4859 ( .B(n1203), .A(n1204), .S(n2553), .Y(n1202) );
  MUX2X1 U4860 ( .B(n1206), .A(n1207), .S(n2553), .Y(n1205) );
  MUX2X1 U4861 ( .B(n1209), .A(n1210), .S(n2553), .Y(n1208) );
  MUX2X1 U4862 ( .B(n1212), .A(n1213), .S(n2628), .Y(n1211) );
  MUX2X1 U4863 ( .B(n1214), .A(n1215), .S(n18), .Y(data_out[13]) );
  MUX2X1 U4864 ( .B(n1217), .A(n1218), .S(n2553), .Y(n1216) );
  MUX2X1 U4865 ( .B(n1220), .A(n1221), .S(n2553), .Y(n1219) );
  MUX2X1 U4866 ( .B(n1223), .A(n1224), .S(n2553), .Y(n1222) );
  MUX2X1 U4867 ( .B(n1226), .A(n1227), .S(n2553), .Y(n1225) );
  MUX2X1 U4868 ( .B(n1229), .A(n1230), .S(n2628), .Y(n1228) );
  MUX2X1 U4869 ( .B(n1232), .A(n1233), .S(n2554), .Y(n1231) );
  MUX2X1 U4870 ( .B(n1235), .A(n1236), .S(n2554), .Y(n1234) );
  MUX2X1 U4871 ( .B(n1238), .A(n1239), .S(n2554), .Y(n1237) );
  MUX2X1 U4872 ( .B(n1241), .A(n1242), .S(n2554), .Y(n1240) );
  MUX2X1 U4873 ( .B(n1244), .A(n1245), .S(n2628), .Y(n1243) );
  MUX2X1 U4874 ( .B(n1247), .A(n1248), .S(n2554), .Y(n1246) );
  MUX2X1 U4875 ( .B(n1250), .A(n1251), .S(n2554), .Y(n1249) );
  MUX2X1 U4876 ( .B(n1253), .A(n1254), .S(n2554), .Y(n1252) );
  MUX2X1 U4877 ( .B(n1256), .A(n1257), .S(n2554), .Y(n1255) );
  MUX2X1 U4878 ( .B(n1259), .A(n1260), .S(n2628), .Y(n1258) );
  MUX2X1 U4879 ( .B(n1262), .A(n1263), .S(n2554), .Y(n1261) );
  MUX2X1 U4880 ( .B(n1265), .A(n1266), .S(n2554), .Y(n1264) );
  MUX2X1 U4881 ( .B(n1268), .A(n1269), .S(n2554), .Y(n1267) );
  MUX2X1 U4882 ( .B(n1271), .A(n1272), .S(n2554), .Y(n1270) );
  MUX2X1 U4883 ( .B(n1274), .A(n1275), .S(n2628), .Y(n1273) );
  MUX2X1 U4884 ( .B(n1276), .A(n1277), .S(n18), .Y(data_out[14]) );
  MUX2X1 U4885 ( .B(n1279), .A(n1280), .S(n2555), .Y(n1278) );
  MUX2X1 U4886 ( .B(n1282), .A(n1283), .S(n2555), .Y(n1281) );
  MUX2X1 U4887 ( .B(n1285), .A(n1286), .S(n2555), .Y(n1284) );
  MUX2X1 U4888 ( .B(n1288), .A(n1289), .S(n2555), .Y(n1287) );
  MUX2X1 U4889 ( .B(n1291), .A(n1292), .S(n2629), .Y(n1290) );
  MUX2X1 U4890 ( .B(n1294), .A(n1295), .S(n2555), .Y(n1293) );
  MUX2X1 U4891 ( .B(n1297), .A(n1298), .S(n2555), .Y(n1296) );
  MUX2X1 U4892 ( .B(n1300), .A(n1301), .S(n2555), .Y(n1299) );
  MUX2X1 U4893 ( .B(n1303), .A(n1304), .S(n2555), .Y(n1302) );
  MUX2X1 U4894 ( .B(n1306), .A(n1307), .S(n2629), .Y(n1305) );
  MUX2X1 U4895 ( .B(n1309), .A(n1310), .S(n2555), .Y(n1308) );
  MUX2X1 U4896 ( .B(n1312), .A(n1313), .S(n2555), .Y(n1311) );
  MUX2X1 U4897 ( .B(n1315), .A(n1316), .S(n2555), .Y(n1314) );
  MUX2X1 U4898 ( .B(n1318), .A(n1319), .S(n2555), .Y(n1317) );
  MUX2X1 U4899 ( .B(n1321), .A(n1322), .S(n2629), .Y(n1320) );
  MUX2X1 U4900 ( .B(n1324), .A(n1325), .S(n2556), .Y(n1323) );
  MUX2X1 U4901 ( .B(n1327), .A(n1328), .S(n2556), .Y(n1326) );
  MUX2X1 U4902 ( .B(n1330), .A(n1331), .S(n2556), .Y(n1329) );
  MUX2X1 U4903 ( .B(n1333), .A(n1334), .S(n2556), .Y(n1332) );
  MUX2X1 U4904 ( .B(n1336), .A(n1337), .S(n2629), .Y(n1335) );
  MUX2X1 U4905 ( .B(n1338), .A(n1339), .S(n18), .Y(data_out[15]) );
  MUX2X1 U4906 ( .B(n1341), .A(n1342), .S(n2556), .Y(n1340) );
  MUX2X1 U4907 ( .B(n1344), .A(n1345), .S(n2556), .Y(n1343) );
  MUX2X1 U4908 ( .B(n1347), .A(n1348), .S(n2556), .Y(n1346) );
  MUX2X1 U4909 ( .B(n1350), .A(n1351), .S(n2556), .Y(n1349) );
  MUX2X1 U4910 ( .B(n1353), .A(n1354), .S(n2629), .Y(n1352) );
  MUX2X1 U4911 ( .B(n1356), .A(n1357), .S(n2556), .Y(n1355) );
  MUX2X1 U4912 ( .B(n1359), .A(n1360), .S(n2556), .Y(n1358) );
  MUX2X1 U4913 ( .B(n1362), .A(n1363), .S(n2556), .Y(n1361) );
  MUX2X1 U4914 ( .B(n1365), .A(n1366), .S(n2556), .Y(n1364) );
  MUX2X1 U4915 ( .B(n1368), .A(n1369), .S(n2629), .Y(n1367) );
  MUX2X1 U4916 ( .B(n1371), .A(n1372), .S(n2557), .Y(n1370) );
  MUX2X1 U4917 ( .B(n1374), .A(n1375), .S(n2557), .Y(n1373) );
  MUX2X1 U4918 ( .B(n1377), .A(n1378), .S(n2557), .Y(n1376) );
  MUX2X1 U4919 ( .B(n1380), .A(n1381), .S(n2557), .Y(n1379) );
  MUX2X1 U4920 ( .B(n1383), .A(n1384), .S(n2629), .Y(n1382) );
  MUX2X1 U4921 ( .B(n1386), .A(n1387), .S(n2557), .Y(n1385) );
  MUX2X1 U4922 ( .B(n1389), .A(n1390), .S(n2557), .Y(n1388) );
  MUX2X1 U4923 ( .B(n1392), .A(n1393), .S(n2557), .Y(n1391) );
  MUX2X1 U4924 ( .B(n1395), .A(n1396), .S(n2557), .Y(n1394) );
  MUX2X1 U4925 ( .B(n1398), .A(n1399), .S(n2629), .Y(n1397) );
  MUX2X1 U4926 ( .B(n1400), .A(n1401), .S(n18), .Y(data_out[16]) );
  MUX2X1 U4927 ( .B(n1403), .A(n1404), .S(n2557), .Y(n1402) );
  MUX2X1 U4928 ( .B(n1406), .A(n1407), .S(n2557), .Y(n1405) );
  MUX2X1 U4929 ( .B(n1409), .A(n1410), .S(n2557), .Y(n1408) );
  MUX2X1 U4930 ( .B(n1412), .A(n1413), .S(n2557), .Y(n1411) );
  MUX2X1 U4931 ( .B(n1415), .A(n1416), .S(n2629), .Y(n1414) );
  MUX2X1 U4932 ( .B(n1418), .A(n1419), .S(n2558), .Y(n1417) );
  MUX2X1 U4933 ( .B(n1421), .A(n1422), .S(n2558), .Y(n1420) );
  MUX2X1 U4934 ( .B(n1424), .A(n1425), .S(n2558), .Y(n1423) );
  MUX2X1 U4935 ( .B(n1427), .A(n1428), .S(n2558), .Y(n1426) );
  MUX2X1 U4936 ( .B(n1430), .A(n1431), .S(n2629), .Y(n1429) );
  MUX2X1 U4937 ( .B(n1433), .A(n1434), .S(n2558), .Y(n1432) );
  MUX2X1 U4938 ( .B(n1436), .A(n1437), .S(n2558), .Y(n1435) );
  MUX2X1 U4939 ( .B(n1439), .A(n1440), .S(n2558), .Y(n1438) );
  MUX2X1 U4940 ( .B(n1442), .A(n1443), .S(n2558), .Y(n1441) );
  MUX2X1 U4941 ( .B(n1445), .A(n1446), .S(n2629), .Y(n1444) );
  MUX2X1 U4942 ( .B(n1448), .A(n1449), .S(n2558), .Y(n1447) );
  MUX2X1 U4943 ( .B(n1451), .A(n1452), .S(n2558), .Y(n1450) );
  MUX2X1 U4944 ( .B(n1454), .A(n1455), .S(n2558), .Y(n1453) );
  MUX2X1 U4945 ( .B(n1457), .A(n1458), .S(n2558), .Y(n1456) );
  MUX2X1 U4946 ( .B(n1460), .A(n1461), .S(n2629), .Y(n1459) );
  MUX2X1 U4947 ( .B(n1462), .A(n1463), .S(n18), .Y(data_out[17]) );
  MUX2X1 U4948 ( .B(n1465), .A(n1466), .S(n2559), .Y(n1464) );
  MUX2X1 U4949 ( .B(n1468), .A(n1469), .S(n2559), .Y(n1467) );
  MUX2X1 U4950 ( .B(n1471), .A(n1472), .S(n2559), .Y(n1470) );
  MUX2X1 U4951 ( .B(n1474), .A(n1475), .S(n2559), .Y(n1473) );
  MUX2X1 U4952 ( .B(n1477), .A(n1478), .S(n2630), .Y(n1476) );
  MUX2X1 U4953 ( .B(n1480), .A(n1481), .S(n2559), .Y(n1479) );
  MUX2X1 U4954 ( .B(n1483), .A(n1484), .S(n2559), .Y(n1482) );
  MUX2X1 U4955 ( .B(n1486), .A(n1487), .S(n2559), .Y(n1485) );
  MUX2X1 U4956 ( .B(n1489), .A(n1490), .S(n2559), .Y(n1488) );
  MUX2X1 U4957 ( .B(n1492), .A(n1493), .S(n2630), .Y(n1491) );
  MUX2X1 U4958 ( .B(n1495), .A(n1496), .S(n2559), .Y(n1494) );
  MUX2X1 U4959 ( .B(n1498), .A(n1499), .S(n2559), .Y(n1497) );
  MUX2X1 U4960 ( .B(n1501), .A(n1502), .S(n2559), .Y(n1500) );
  MUX2X1 U4961 ( .B(n1504), .A(n1505), .S(n2559), .Y(n1503) );
  MUX2X1 U4962 ( .B(n1507), .A(n1508), .S(n2630), .Y(n1506) );
  MUX2X1 U4963 ( .B(n1510), .A(n1511), .S(n2560), .Y(n1509) );
  MUX2X1 U4964 ( .B(n1513), .A(n1514), .S(n2560), .Y(n1512) );
  MUX2X1 U4965 ( .B(n1516), .A(n1517), .S(n2560), .Y(n1515) );
  MUX2X1 U4966 ( .B(n1519), .A(n1520), .S(n2560), .Y(n1518) );
  MUX2X1 U4967 ( .B(n1522), .A(n1523), .S(n2630), .Y(n1521) );
  MUX2X1 U4968 ( .B(n1524), .A(n1525), .S(n18), .Y(data_out[18]) );
  MUX2X1 U4969 ( .B(n1527), .A(n1528), .S(n2560), .Y(n1526) );
  MUX2X1 U4970 ( .B(n1530), .A(n1531), .S(n2560), .Y(n1529) );
  MUX2X1 U4971 ( .B(n1533), .A(n1534), .S(n2560), .Y(n1532) );
  MUX2X1 U4972 ( .B(n1536), .A(n1537), .S(n2560), .Y(n1535) );
  MUX2X1 U4973 ( .B(n1539), .A(n1540), .S(n2630), .Y(n1538) );
  MUX2X1 U4974 ( .B(n1542), .A(n1543), .S(n2560), .Y(n1541) );
  MUX2X1 U4975 ( .B(n1545), .A(n1546), .S(n2560), .Y(n1544) );
  MUX2X1 U4976 ( .B(n1548), .A(n1549), .S(n2560), .Y(n1547) );
  MUX2X1 U4977 ( .B(n1551), .A(n1552), .S(n2560), .Y(n1550) );
  MUX2X1 U4978 ( .B(n1554), .A(n1555), .S(n2630), .Y(n1553) );
  MUX2X1 U4979 ( .B(n1557), .A(n1558), .S(n2561), .Y(n1556) );
  MUX2X1 U4980 ( .B(n1560), .A(n1561), .S(n2561), .Y(n1559) );
  MUX2X1 U4981 ( .B(n1563), .A(n1564), .S(n2561), .Y(n1562) );
  MUX2X1 U4982 ( .B(n1566), .A(n1567), .S(n2561), .Y(n1565) );
  MUX2X1 U4983 ( .B(n1569), .A(n1570), .S(n2630), .Y(n1568) );
  MUX2X1 U4984 ( .B(n1572), .A(n1573), .S(n2561), .Y(n1571) );
  MUX2X1 U4985 ( .B(n1575), .A(n1576), .S(n2561), .Y(n1574) );
  MUX2X1 U4986 ( .B(n1578), .A(n1579), .S(n2561), .Y(n1577) );
  MUX2X1 U4987 ( .B(n1581), .A(n1582), .S(n2561), .Y(n1580) );
  MUX2X1 U4988 ( .B(n1584), .A(n1585), .S(n2630), .Y(n1583) );
  MUX2X1 U4989 ( .B(n1586), .A(n1587), .S(n18), .Y(data_out[19]) );
  MUX2X1 U4990 ( .B(n1589), .A(n1590), .S(n2561), .Y(n1588) );
  MUX2X1 U4991 ( .B(n1592), .A(n1593), .S(n2561), .Y(n1591) );
  MUX2X1 U4992 ( .B(n1595), .A(n1596), .S(n2561), .Y(n1594) );
  MUX2X1 U4993 ( .B(n1598), .A(n1599), .S(n2561), .Y(n1597) );
  MUX2X1 U4994 ( .B(n1601), .A(n1602), .S(n2630), .Y(n1600) );
  MUX2X1 U4995 ( .B(n1604), .A(n1605), .S(n2562), .Y(n1603) );
  MUX2X1 U4996 ( .B(n1607), .A(n1608), .S(n2562), .Y(n1606) );
  MUX2X1 U4997 ( .B(n1610), .A(n1611), .S(n2562), .Y(n1609) );
  MUX2X1 U4998 ( .B(n1613), .A(n1614), .S(n2562), .Y(n1612) );
  MUX2X1 U4999 ( .B(n1616), .A(n1617), .S(n2630), .Y(n1615) );
  MUX2X1 U5000 ( .B(n1619), .A(n1620), .S(n2562), .Y(n1618) );
  MUX2X1 U5001 ( .B(n1622), .A(n1623), .S(n2562), .Y(n1621) );
  MUX2X1 U5002 ( .B(n1625), .A(n1626), .S(n2562), .Y(n1624) );
  MUX2X1 U5003 ( .B(n1628), .A(n1629), .S(n2562), .Y(n1627) );
  MUX2X1 U5004 ( .B(n1631), .A(n1632), .S(n2630), .Y(n1630) );
  MUX2X1 U5005 ( .B(n1634), .A(n1635), .S(n2562), .Y(n1633) );
  MUX2X1 U5006 ( .B(n1637), .A(n1638), .S(n2562), .Y(n1636) );
  MUX2X1 U5007 ( .B(n1640), .A(n1641), .S(n2562), .Y(n1639) );
  MUX2X1 U5008 ( .B(n1643), .A(n1644), .S(n2562), .Y(n1642) );
  MUX2X1 U5009 ( .B(n1646), .A(n1647), .S(n2630), .Y(n1645) );
  MUX2X1 U5010 ( .B(n1648), .A(n1649), .S(n18), .Y(data_out[20]) );
  MUX2X1 U5011 ( .B(n1651), .A(n1652), .S(n2563), .Y(n1650) );
  MUX2X1 U5012 ( .B(n1654), .A(n1655), .S(n2563), .Y(n1653) );
  MUX2X1 U5013 ( .B(n1657), .A(n1658), .S(n2563), .Y(n1656) );
  MUX2X1 U5014 ( .B(n1660), .A(n1661), .S(n2563), .Y(n1659) );
  MUX2X1 U5015 ( .B(n1663), .A(n1664), .S(n2631), .Y(n1662) );
  MUX2X1 U5016 ( .B(n1666), .A(n1667), .S(n2563), .Y(n1665) );
  MUX2X1 U5017 ( .B(n1669), .A(n1670), .S(n2563), .Y(n1668) );
  MUX2X1 U5018 ( .B(n1672), .A(n1673), .S(n2563), .Y(n1671) );
  MUX2X1 U5019 ( .B(n1675), .A(n1676), .S(n2563), .Y(n1674) );
  MUX2X1 U5020 ( .B(n1678), .A(n1679), .S(n2631), .Y(n1677) );
  MUX2X1 U5021 ( .B(n1681), .A(n1682), .S(n2563), .Y(n1680) );
  MUX2X1 U5022 ( .B(n1684), .A(n1685), .S(n2563), .Y(n1683) );
  MUX2X1 U5023 ( .B(n1687), .A(n1688), .S(n2563), .Y(n1686) );
  MUX2X1 U5024 ( .B(n1690), .A(n1691), .S(n2563), .Y(n1689) );
  MUX2X1 U5025 ( .B(n1693), .A(n1694), .S(n2631), .Y(n1692) );
  MUX2X1 U5026 ( .B(n1696), .A(n1697), .S(n2564), .Y(n1695) );
  MUX2X1 U5027 ( .B(n1699), .A(n1700), .S(n2564), .Y(n1698) );
  MUX2X1 U5028 ( .B(n1702), .A(n1703), .S(n2564), .Y(n1701) );
  MUX2X1 U5029 ( .B(n1705), .A(n1706), .S(n2564), .Y(n1704) );
  MUX2X1 U5030 ( .B(n1708), .A(n1709), .S(n2631), .Y(n1707) );
  MUX2X1 U5031 ( .B(n1710), .A(n1711), .S(n18), .Y(data_out[21]) );
  MUX2X1 U5032 ( .B(n1713), .A(n1714), .S(n2564), .Y(n1712) );
  MUX2X1 U5033 ( .B(n1716), .A(n1717), .S(n2564), .Y(n1715) );
  MUX2X1 U5034 ( .B(n1719), .A(n1720), .S(n2564), .Y(n1718) );
  MUX2X1 U5035 ( .B(n1722), .A(n1723), .S(n2564), .Y(n1721) );
  MUX2X1 U5036 ( .B(n1725), .A(n1726), .S(n2631), .Y(n1724) );
  MUX2X1 U5037 ( .B(n1728), .A(n1729), .S(n2564), .Y(n1727) );
  MUX2X1 U5038 ( .B(n1731), .A(n1732), .S(n2564), .Y(n1730) );
  MUX2X1 U5039 ( .B(n1734), .A(n1735), .S(n2564), .Y(n1733) );
  MUX2X1 U5040 ( .B(n1737), .A(n1738), .S(n2564), .Y(n1736) );
  MUX2X1 U5041 ( .B(n1740), .A(n1741), .S(n2631), .Y(n1739) );
  MUX2X1 U5042 ( .B(n1743), .A(n1744), .S(n2565), .Y(n1742) );
  MUX2X1 U5043 ( .B(n1746), .A(n1747), .S(n2565), .Y(n1745) );
  MUX2X1 U5044 ( .B(n1749), .A(n1750), .S(n2565), .Y(n1748) );
  MUX2X1 U5045 ( .B(n1752), .A(n1753), .S(n2565), .Y(n1751) );
  MUX2X1 U5046 ( .B(n1755), .A(n1756), .S(n2631), .Y(n1754) );
  MUX2X1 U5047 ( .B(n1758), .A(n1759), .S(n2565), .Y(n1757) );
  MUX2X1 U5048 ( .B(n1761), .A(n1762), .S(n2565), .Y(n1760) );
  MUX2X1 U5049 ( .B(n1764), .A(n1765), .S(n2565), .Y(n1763) );
  MUX2X1 U5050 ( .B(n1767), .A(n1768), .S(n2565), .Y(n1766) );
  MUX2X1 U5051 ( .B(n1770), .A(n1771), .S(n2631), .Y(n1769) );
  MUX2X1 U5052 ( .B(n1772), .A(n1773), .S(n18), .Y(data_out[22]) );
  MUX2X1 U5053 ( .B(n1775), .A(n1776), .S(n2565), .Y(n1774) );
  MUX2X1 U5054 ( .B(n1778), .A(n1779), .S(n2565), .Y(n1777) );
  MUX2X1 U5055 ( .B(n1781), .A(n1782), .S(n2565), .Y(n1780) );
  MUX2X1 U5056 ( .B(n1784), .A(n1785), .S(n2565), .Y(n1783) );
  MUX2X1 U5057 ( .B(n1787), .A(n1788), .S(n2631), .Y(n1786) );
  MUX2X1 U5058 ( .B(n1790), .A(n1791), .S(n2566), .Y(n1789) );
  MUX2X1 U5059 ( .B(n1793), .A(n1794), .S(n2566), .Y(n1792) );
  MUX2X1 U5060 ( .B(n1796), .A(n1797), .S(n2566), .Y(n1795) );
  MUX2X1 U5061 ( .B(n1799), .A(n1800), .S(n2566), .Y(n1798) );
  MUX2X1 U5062 ( .B(n1802), .A(n1803), .S(n2631), .Y(n1801) );
  MUX2X1 U5063 ( .B(n1805), .A(n1806), .S(n2566), .Y(n1804) );
  MUX2X1 U5064 ( .B(n1808), .A(n1809), .S(n2566), .Y(n1807) );
  MUX2X1 U5065 ( .B(n1811), .A(n1812), .S(n2566), .Y(n1810) );
  MUX2X1 U5066 ( .B(n1814), .A(n1815), .S(n2566), .Y(n1813) );
  MUX2X1 U5067 ( .B(n1817), .A(n1818), .S(n2631), .Y(n1816) );
  MUX2X1 U5068 ( .B(n1820), .A(n1821), .S(n2566), .Y(n1819) );
  MUX2X1 U5069 ( .B(n1823), .A(n1824), .S(n2566), .Y(n1822) );
  MUX2X1 U5070 ( .B(n1826), .A(n1827), .S(n2566), .Y(n1825) );
  MUX2X1 U5071 ( .B(n1829), .A(n1830), .S(n2566), .Y(n1828) );
  MUX2X1 U5072 ( .B(n1832), .A(n1833), .S(n2631), .Y(n1831) );
  MUX2X1 U5073 ( .B(n1834), .A(n1835), .S(n18), .Y(data_out[23]) );
  MUX2X1 U5074 ( .B(n1837), .A(n1838), .S(n2567), .Y(n1836) );
  MUX2X1 U5075 ( .B(n1840), .A(n1841), .S(n2567), .Y(n1839) );
  MUX2X1 U5076 ( .B(n1843), .A(n1844), .S(n2567), .Y(n1842) );
  MUX2X1 U5077 ( .B(n1846), .A(n1847), .S(n2567), .Y(n1845) );
  MUX2X1 U5078 ( .B(n1849), .A(n1850), .S(n2632), .Y(n1848) );
  MUX2X1 U5079 ( .B(n1852), .A(n1853), .S(n2567), .Y(n1851) );
  MUX2X1 U5080 ( .B(n1855), .A(n1856), .S(n2567), .Y(n1854) );
  MUX2X1 U5081 ( .B(n1858), .A(n1859), .S(n2567), .Y(n1857) );
  MUX2X1 U5082 ( .B(n1861), .A(n1862), .S(n2567), .Y(n1860) );
  MUX2X1 U5083 ( .B(n1864), .A(n1865), .S(n2632), .Y(n1863) );
  MUX2X1 U5084 ( .B(n1867), .A(n1868), .S(n2567), .Y(n1866) );
  MUX2X1 U5085 ( .B(n1870), .A(n1871), .S(n2567), .Y(n1869) );
  MUX2X1 U5086 ( .B(n1873), .A(n1874), .S(n2567), .Y(n1872) );
  MUX2X1 U5087 ( .B(n1876), .A(n1877), .S(n2567), .Y(n1875) );
  MUX2X1 U5088 ( .B(n1879), .A(n1880), .S(n2632), .Y(n1878) );
  MUX2X1 U5089 ( .B(n1882), .A(n1883), .S(n2568), .Y(n1881) );
  MUX2X1 U5090 ( .B(n1885), .A(n1886), .S(n2568), .Y(n1884) );
  MUX2X1 U5091 ( .B(n1888), .A(n1889), .S(n2568), .Y(n1887) );
  MUX2X1 U5092 ( .B(n1891), .A(n1892), .S(n2568), .Y(n1890) );
  MUX2X1 U5093 ( .B(n1894), .A(n1895), .S(n2632), .Y(n1893) );
  MUX2X1 U5094 ( .B(n1896), .A(n1897), .S(n18), .Y(data_out[24]) );
  MUX2X1 U5095 ( .B(n1899), .A(n1900), .S(n2568), .Y(n1898) );
  MUX2X1 U5096 ( .B(n1902), .A(n1903), .S(n2568), .Y(n1901) );
  MUX2X1 U5097 ( .B(n1905), .A(n1906), .S(n2568), .Y(n1904) );
  MUX2X1 U5098 ( .B(n1908), .A(n1909), .S(n2568), .Y(n1907) );
  MUX2X1 U5099 ( .B(n1911), .A(n1912), .S(n2632), .Y(n1910) );
  MUX2X1 U5100 ( .B(n1914), .A(n1915), .S(n2568), .Y(n1913) );
  MUX2X1 U5101 ( .B(n1917), .A(n1918), .S(n2568), .Y(n1916) );
  MUX2X1 U5102 ( .B(n1920), .A(n1921), .S(n2568), .Y(n1919) );
  MUX2X1 U5103 ( .B(n1923), .A(n1924), .S(n2568), .Y(n1922) );
  MUX2X1 U5104 ( .B(n1926), .A(n1927), .S(n2632), .Y(n1925) );
  MUX2X1 U5105 ( .B(n1929), .A(n1930), .S(n2569), .Y(n1928) );
  MUX2X1 U5106 ( .B(n1932), .A(n1933), .S(n2569), .Y(n1931) );
  MUX2X1 U5107 ( .B(n1935), .A(n1936), .S(n2569), .Y(n1934) );
  MUX2X1 U5108 ( .B(n1938), .A(n1939), .S(n2569), .Y(n1937) );
  MUX2X1 U5109 ( .B(n1941), .A(n1942), .S(n2632), .Y(n1940) );
  MUX2X1 U5110 ( .B(n1944), .A(n1945), .S(n2569), .Y(n1943) );
  MUX2X1 U5111 ( .B(n1947), .A(n1948), .S(n2569), .Y(n1946) );
  MUX2X1 U5112 ( .B(n1950), .A(n1951), .S(n2569), .Y(n1949) );
  MUX2X1 U5113 ( .B(n1953), .A(n1954), .S(n2569), .Y(n1952) );
  MUX2X1 U5114 ( .B(n1956), .A(n1957), .S(n2632), .Y(n1955) );
  MUX2X1 U5115 ( .B(n1958), .A(n1959), .S(n18), .Y(data_out[25]) );
  MUX2X1 U5116 ( .B(n1961), .A(n1962), .S(n2569), .Y(n1960) );
  MUX2X1 U5117 ( .B(n1964), .A(n1965), .S(n2569), .Y(n1963) );
  MUX2X1 U5118 ( .B(n1967), .A(n1968), .S(n2569), .Y(n1966) );
  MUX2X1 U5119 ( .B(n1970), .A(n1971), .S(n2569), .Y(n1969) );
  MUX2X1 U5120 ( .B(n1973), .A(n1974), .S(n2632), .Y(n1972) );
  MUX2X1 U5121 ( .B(n1976), .A(n1977), .S(n2570), .Y(n1975) );
  MUX2X1 U5122 ( .B(n1979), .A(n1980), .S(n2570), .Y(n1978) );
  MUX2X1 U5123 ( .B(n1982), .A(n1983), .S(n2570), .Y(n1981) );
  MUX2X1 U5124 ( .B(n1985), .A(n1986), .S(n2570), .Y(n1984) );
  MUX2X1 U5125 ( .B(n1988), .A(n1989), .S(n2632), .Y(n1987) );
  MUX2X1 U5126 ( .B(n1991), .A(n1992), .S(n2570), .Y(n1990) );
  MUX2X1 U5127 ( .B(n1994), .A(n1995), .S(n2570), .Y(n1993) );
  MUX2X1 U5128 ( .B(n1997), .A(n1998), .S(n2570), .Y(n1996) );
  MUX2X1 U5129 ( .B(n2000), .A(n2001), .S(n2570), .Y(n1999) );
  MUX2X1 U5130 ( .B(n2003), .A(n2004), .S(n2632), .Y(n2002) );
  MUX2X1 U5131 ( .B(n2006), .A(n2007), .S(n2570), .Y(n2005) );
  MUX2X1 U5132 ( .B(n2009), .A(n2010), .S(n2570), .Y(n2008) );
  MUX2X1 U5133 ( .B(n2012), .A(n2013), .S(n2570), .Y(n2011) );
  MUX2X1 U5134 ( .B(n2015), .A(n2016), .S(n2570), .Y(n2014) );
  MUX2X1 U5135 ( .B(n2018), .A(n2019), .S(n2632), .Y(n2017) );
  MUX2X1 U5136 ( .B(n2020), .A(n2021), .S(n18), .Y(data_out[26]) );
  MUX2X1 U5137 ( .B(n2023), .A(n2024), .S(n2571), .Y(n2022) );
  MUX2X1 U5138 ( .B(n2026), .A(n2027), .S(n2571), .Y(n2025) );
  MUX2X1 U5139 ( .B(n2029), .A(n2030), .S(n2571), .Y(n2028) );
  MUX2X1 U5140 ( .B(n2032), .A(n2033), .S(n2571), .Y(n2031) );
  MUX2X1 U5141 ( .B(n2035), .A(n2036), .S(n2633), .Y(n2034) );
  MUX2X1 U5142 ( .B(n2038), .A(n2039), .S(n2571), .Y(n2037) );
  MUX2X1 U5143 ( .B(n2041), .A(n2042), .S(n2571), .Y(n2040) );
  MUX2X1 U5144 ( .B(n2044), .A(n2045), .S(n2571), .Y(n2043) );
  MUX2X1 U5145 ( .B(n2047), .A(n2048), .S(n2571), .Y(n2046) );
  MUX2X1 U5146 ( .B(n2050), .A(n2051), .S(n2633), .Y(n2049) );
  MUX2X1 U5147 ( .B(n2053), .A(n2054), .S(n2571), .Y(n2052) );
  MUX2X1 U5148 ( .B(n2056), .A(n2057), .S(n2571), .Y(n2055) );
  MUX2X1 U5149 ( .B(n2059), .A(n2060), .S(n2571), .Y(n2058) );
  MUX2X1 U5150 ( .B(n2062), .A(n2063), .S(n2571), .Y(n2061) );
  MUX2X1 U5151 ( .B(n2065), .A(n2066), .S(n2633), .Y(n2064) );
  MUX2X1 U5152 ( .B(n2068), .A(n2069), .S(n2572), .Y(n2067) );
  MUX2X1 U5153 ( .B(n2071), .A(n2072), .S(n2572), .Y(n2070) );
  MUX2X1 U5154 ( .B(n2074), .A(n2075), .S(n2572), .Y(n2073) );
  MUX2X1 U5155 ( .B(n2077), .A(n2078), .S(n2572), .Y(n2076) );
  MUX2X1 U5156 ( .B(n2080), .A(n2081), .S(n2633), .Y(n2079) );
  MUX2X1 U5157 ( .B(n2082), .A(n2083), .S(n18), .Y(data_out[27]) );
  MUX2X1 U5158 ( .B(n2085), .A(n2086), .S(n2572), .Y(n2084) );
  MUX2X1 U5159 ( .B(n2088), .A(n2089), .S(n2572), .Y(n2087) );
  MUX2X1 U5160 ( .B(n2091), .A(n2092), .S(n2572), .Y(n2090) );
  MUX2X1 U5161 ( .B(n2094), .A(n2095), .S(n2572), .Y(n2093) );
  MUX2X1 U5162 ( .B(n2097), .A(n2098), .S(n2633), .Y(n2096) );
  MUX2X1 U5163 ( .B(n2100), .A(n2101), .S(n2572), .Y(n2099) );
  MUX2X1 U5164 ( .B(n2103), .A(n2104), .S(n2572), .Y(n2102) );
  MUX2X1 U5165 ( .B(n2106), .A(n2107), .S(n2572), .Y(n2105) );
  MUX2X1 U5166 ( .B(n2109), .A(n2110), .S(n2572), .Y(n2108) );
  MUX2X1 U5167 ( .B(n2112), .A(n2113), .S(n2633), .Y(n2111) );
  MUX2X1 U5168 ( .B(n2115), .A(n2116), .S(n2573), .Y(n2114) );
  MUX2X1 U5169 ( .B(n2118), .A(n2119), .S(n2573), .Y(n2117) );
  MUX2X1 U5170 ( .B(n2121), .A(n2122), .S(n2573), .Y(n2120) );
  MUX2X1 U5171 ( .B(n2124), .A(n2125), .S(n2573), .Y(n2123) );
  MUX2X1 U5172 ( .B(n2127), .A(n2128), .S(n2633), .Y(n2126) );
  MUX2X1 U5173 ( .B(n2130), .A(n2131), .S(n2573), .Y(n2129) );
  MUX2X1 U5174 ( .B(n2133), .A(n2134), .S(n2573), .Y(n2132) );
  MUX2X1 U5175 ( .B(n2136), .A(n2137), .S(n2573), .Y(n2135) );
  MUX2X1 U5176 ( .B(n2139), .A(n2140), .S(n2573), .Y(n2138) );
  MUX2X1 U5177 ( .B(n2142), .A(n2143), .S(n2633), .Y(n2141) );
  MUX2X1 U5178 ( .B(n2144), .A(n2145), .S(n18), .Y(data_out[28]) );
  MUX2X1 U5179 ( .B(n2147), .A(n2148), .S(n2573), .Y(n2146) );
  MUX2X1 U5180 ( .B(n2150), .A(n2151), .S(n2573), .Y(n2149) );
  MUX2X1 U5181 ( .B(n2153), .A(n2154), .S(n2573), .Y(n2152) );
  MUX2X1 U5182 ( .B(n2156), .A(n2157), .S(n2573), .Y(n2155) );
  MUX2X1 U5183 ( .B(n2159), .A(n2160), .S(n2633), .Y(n2158) );
  MUX2X1 U5184 ( .B(n2162), .A(n2163), .S(n2574), .Y(n2161) );
  MUX2X1 U5185 ( .B(n2165), .A(n2166), .S(n2574), .Y(n2164) );
  MUX2X1 U5186 ( .B(n2168), .A(n2169), .S(n2574), .Y(n2167) );
  MUX2X1 U5187 ( .B(n2171), .A(n2172), .S(n2574), .Y(n2170) );
  MUX2X1 U5188 ( .B(n2174), .A(n2175), .S(n2633), .Y(n2173) );
  MUX2X1 U5189 ( .B(n2177), .A(n2178), .S(n2574), .Y(n2176) );
  MUX2X1 U5190 ( .B(n2180), .A(n2181), .S(n2574), .Y(n2179) );
  MUX2X1 U5191 ( .B(n2183), .A(n2184), .S(n2574), .Y(n2182) );
  MUX2X1 U5192 ( .B(n2186), .A(n2187), .S(n2574), .Y(n2185) );
  MUX2X1 U5193 ( .B(n2189), .A(n2190), .S(n2633), .Y(n2188) );
  MUX2X1 U5194 ( .B(n2192), .A(n2193), .S(n2574), .Y(n2191) );
  MUX2X1 U5195 ( .B(n2195), .A(n2196), .S(n2574), .Y(n2194) );
  MUX2X1 U5196 ( .B(n2198), .A(n2199), .S(n2574), .Y(n2197) );
  MUX2X1 U5197 ( .B(n2201), .A(n2202), .S(n2574), .Y(n2200) );
  MUX2X1 U5198 ( .B(n2204), .A(n2205), .S(n2633), .Y(n2203) );
  MUX2X1 U5199 ( .B(n2206), .A(n2207), .S(n18), .Y(data_out[29]) );
  MUX2X1 U5200 ( .B(n2209), .A(n2210), .S(n2575), .Y(n2208) );
  MUX2X1 U5201 ( .B(n2212), .A(n2226), .S(n2575), .Y(n2211) );
  MUX2X1 U5202 ( .B(n2228), .A(n2229), .S(n2575), .Y(n2227) );
  MUX2X1 U5203 ( .B(n2231), .A(n2232), .S(n2575), .Y(n2230) );
  MUX2X1 U5204 ( .B(n2234), .A(n2235), .S(n2634), .Y(n2233) );
  MUX2X1 U5205 ( .B(n2237), .A(n2238), .S(n2575), .Y(n2236) );
  MUX2X1 U5206 ( .B(n2240), .A(n2241), .S(n2575), .Y(n2239) );
  MUX2X1 U5207 ( .B(n2243), .A(n2244), .S(n2575), .Y(n2242) );
  MUX2X1 U5208 ( .B(n2246), .A(n2247), .S(n2575), .Y(n2245) );
  MUX2X1 U5209 ( .B(n2249), .A(n2250), .S(n2634), .Y(n2248) );
  MUX2X1 U5210 ( .B(n2252), .A(n2253), .S(n2575), .Y(n2251) );
  MUX2X1 U5211 ( .B(n2255), .A(n2256), .S(n2575), .Y(n2254) );
  MUX2X1 U5212 ( .B(n2258), .A(n2259), .S(n2575), .Y(n2257) );
  MUX2X1 U5213 ( .B(n2261), .A(n2262), .S(n2575), .Y(n2260) );
  MUX2X1 U5214 ( .B(n2264), .A(n2265), .S(n2634), .Y(n2263) );
  MUX2X1 U5215 ( .B(n2267), .A(n2268), .S(n2576), .Y(n2266) );
  MUX2X1 U5216 ( .B(n2270), .A(n2271), .S(n2576), .Y(n2269) );
  MUX2X1 U5217 ( .B(n2273), .A(n2274), .S(n2576), .Y(n2272) );
  MUX2X1 U5218 ( .B(n2276), .A(n2277), .S(n2576), .Y(n2275) );
  MUX2X1 U5219 ( .B(n2279), .A(n2280), .S(n2634), .Y(n2278) );
  MUX2X1 U5220 ( .B(n2281), .A(n2282), .S(n18), .Y(data_out[30]) );
  MUX2X1 U5221 ( .B(n2284), .A(n2285), .S(n2576), .Y(n2283) );
  MUX2X1 U5222 ( .B(n2287), .A(n2288), .S(n2576), .Y(n2286) );
  MUX2X1 U5223 ( .B(n2290), .A(n2291), .S(n2576), .Y(n2289) );
  MUX2X1 U5224 ( .B(n2293), .A(n2294), .S(n2576), .Y(n2292) );
  MUX2X1 U5225 ( .B(n2296), .A(n2297), .S(n2634), .Y(n2295) );
  MUX2X1 U5226 ( .B(n2299), .A(n2300), .S(n2576), .Y(n2298) );
  MUX2X1 U5227 ( .B(n2302), .A(n2303), .S(n2576), .Y(n2301) );
  MUX2X1 U5228 ( .B(n2305), .A(n2306), .S(n2576), .Y(n2304) );
  MUX2X1 U5229 ( .B(n2308), .A(n2309), .S(n2576), .Y(n2307) );
  MUX2X1 U5230 ( .B(n2311), .A(n2312), .S(n2634), .Y(n2310) );
  MUX2X1 U5231 ( .B(n2314), .A(n2315), .S(n2577), .Y(n2313) );
  MUX2X1 U5232 ( .B(n2317), .A(n2318), .S(n2577), .Y(n2316) );
  MUX2X1 U5233 ( .B(n2320), .A(n2321), .S(n2577), .Y(n2319) );
  MUX2X1 U5234 ( .B(n2323), .A(n2324), .S(n2577), .Y(n2322) );
  MUX2X1 U5235 ( .B(n2326), .A(n2327), .S(n2634), .Y(n2325) );
  MUX2X1 U5236 ( .B(n2329), .A(n2330), .S(n2577), .Y(n2328) );
  MUX2X1 U5237 ( .B(n2332), .A(n2333), .S(n2577), .Y(n2331) );
  MUX2X1 U5238 ( .B(n2335), .A(n2336), .S(n2577), .Y(n2334) );
  MUX2X1 U5239 ( .B(n2338), .A(n2339), .S(n2577), .Y(n2337) );
  MUX2X1 U5240 ( .B(n2341), .A(n2342), .S(n2634), .Y(n2340) );
  MUX2X1 U5241 ( .B(n2343), .A(n2344), .S(n18), .Y(data_out[31]) );
  MUX2X1 U5242 ( .B(n2346), .A(n2347), .S(n2577), .Y(n2345) );
  MUX2X1 U5243 ( .B(n2349), .A(n2350), .S(n2577), .Y(n2348) );
  MUX2X1 U5244 ( .B(n2352), .A(n2353), .S(n2577), .Y(n2351) );
  MUX2X1 U5245 ( .B(n2355), .A(n2356), .S(n2577), .Y(n2354) );
  MUX2X1 U5246 ( .B(n2358), .A(n2359), .S(n2634), .Y(n2357) );
  MUX2X1 U5247 ( .B(n2361), .A(n2362), .S(n2578), .Y(n2360) );
  MUX2X1 U5248 ( .B(n2364), .A(n2365), .S(n2578), .Y(n2363) );
  MUX2X1 U5249 ( .B(n2367), .A(n2368), .S(n2578), .Y(n2366) );
  MUX2X1 U5250 ( .B(n2370), .A(n2371), .S(n2578), .Y(n2369) );
  MUX2X1 U5251 ( .B(n2373), .A(n2374), .S(n2634), .Y(n2372) );
  MUX2X1 U5252 ( .B(n2376), .A(n2377), .S(n2578), .Y(n2375) );
  MUX2X1 U5253 ( .B(n2379), .A(n2380), .S(n2578), .Y(n2378) );
  MUX2X1 U5254 ( .B(n2382), .A(n2383), .S(n2578), .Y(n2381) );
  MUX2X1 U5255 ( .B(n2385), .A(n2386), .S(n2578), .Y(n2384) );
  MUX2X1 U5256 ( .B(n2388), .A(n2389), .S(n2634), .Y(n2387) );
  MUX2X1 U5257 ( .B(n2391), .A(n2392), .S(n2578), .Y(n2390) );
  MUX2X1 U5258 ( .B(n2394), .A(n2395), .S(n2578), .Y(n2393) );
  MUX2X1 U5259 ( .B(n2397), .A(n2398), .S(n2578), .Y(n2396) );
  MUX2X1 U5260 ( .B(n2400), .A(n2401), .S(n2578), .Y(n2399) );
  MUX2X1 U5261 ( .B(n2403), .A(n2404), .S(n2634), .Y(n2402) );
  MUX2X1 U5262 ( .B(n2405), .A(n2406), .S(n18), .Y(data_out[32]) );
  MUX2X1 U5263 ( .B(arr[2046]), .A(arr[2079]), .S(n2437), .Y(n350) );
  MUX2X1 U5264 ( .B(arr[1980]), .A(arr[2013]), .S(n2437), .Y(n349) );
  MUX2X1 U5265 ( .B(arr[1914]), .A(arr[1947]), .S(n2437), .Y(n353) );
  MUX2X1 U5266 ( .B(arr[1848]), .A(arr[1881]), .S(n2437), .Y(n352) );
  MUX2X1 U5267 ( .B(n351), .A(n348), .S(n2594), .Y(n362) );
  MUX2X1 U5268 ( .B(arr[1782]), .A(arr[1815]), .S(n2437), .Y(n356) );
  MUX2X1 U5269 ( .B(arr[1716]), .A(arr[1749]), .S(n2437), .Y(n355) );
  MUX2X1 U5270 ( .B(arr[1650]), .A(arr[1683]), .S(n2437), .Y(n359) );
  MUX2X1 U5271 ( .B(arr[1584]), .A(arr[1617]), .S(n2437), .Y(n358) );
  MUX2X1 U5272 ( .B(n357), .A(n354), .S(n2594), .Y(n361) );
  MUX2X1 U5273 ( .B(arr[1518]), .A(arr[1551]), .S(n2437), .Y(n365) );
  MUX2X1 U5274 ( .B(arr[1452]), .A(arr[1485]), .S(n2437), .Y(n364) );
  MUX2X1 U5275 ( .B(arr[1386]), .A(arr[1419]), .S(n2437), .Y(n368) );
  MUX2X1 U5276 ( .B(arr[1320]), .A(arr[1353]), .S(n2437), .Y(n367) );
  MUX2X1 U5277 ( .B(n366), .A(n363), .S(n2594), .Y(n377) );
  MUX2X1 U5278 ( .B(arr[1254]), .A(arr[1287]), .S(n2438), .Y(n371) );
  MUX2X1 U5279 ( .B(arr[1188]), .A(arr[1221]), .S(n2438), .Y(n370) );
  MUX2X1 U5280 ( .B(arr[1122]), .A(arr[1155]), .S(n2438), .Y(n374) );
  MUX2X1 U5281 ( .B(arr[1056]), .A(arr[1089]), .S(n2438), .Y(n373) );
  MUX2X1 U5282 ( .B(n372), .A(n369), .S(n2594), .Y(n376) );
  MUX2X1 U5283 ( .B(n375), .A(n360), .S(n2635), .Y(n409) );
  MUX2X1 U5284 ( .B(arr[990]), .A(arr[1023]), .S(n2438), .Y(n380) );
  MUX2X1 U5285 ( .B(arr[924]), .A(arr[957]), .S(n2438), .Y(n379) );
  MUX2X1 U5286 ( .B(arr[858]), .A(arr[891]), .S(n2438), .Y(n383) );
  MUX2X1 U5287 ( .B(arr[792]), .A(arr[825]), .S(n2438), .Y(n382) );
  MUX2X1 U5288 ( .B(n381), .A(n378), .S(n2594), .Y(n392) );
  MUX2X1 U5289 ( .B(arr[726]), .A(arr[759]), .S(n2438), .Y(n386) );
  MUX2X1 U5290 ( .B(arr[660]), .A(arr[693]), .S(n2438), .Y(n385) );
  MUX2X1 U5291 ( .B(arr[594]), .A(arr[627]), .S(n2438), .Y(n389) );
  MUX2X1 U5292 ( .B(arr[528]), .A(arr[561]), .S(n2438), .Y(n388) );
  MUX2X1 U5293 ( .B(n387), .A(n384), .S(n2594), .Y(n391) );
  MUX2X1 U5294 ( .B(arr[462]), .A(arr[495]), .S(n2439), .Y(n395) );
  MUX2X1 U5295 ( .B(arr[396]), .A(arr[429]), .S(n2439), .Y(n394) );
  MUX2X1 U5296 ( .B(arr[330]), .A(arr[363]), .S(n2439), .Y(n398) );
  MUX2X1 U5297 ( .B(arr[264]), .A(arr[297]), .S(n2439), .Y(n397) );
  MUX2X1 U5298 ( .B(n396), .A(n393), .S(n2594), .Y(n407) );
  MUX2X1 U5299 ( .B(arr[198]), .A(arr[231]), .S(n2439), .Y(n401) );
  MUX2X1 U5300 ( .B(arr[132]), .A(arr[165]), .S(n2439), .Y(n400) );
  MUX2X1 U5301 ( .B(arr[66]), .A(arr[99]), .S(n2439), .Y(n404) );
  MUX2X1 U5302 ( .B(arr[0]), .A(arr[33]), .S(n2439), .Y(n403) );
  MUX2X1 U5303 ( .B(n402), .A(n399), .S(n2594), .Y(n406) );
  MUX2X1 U5304 ( .B(n405), .A(n390), .S(n2635), .Y(n408) );
  MUX2X1 U5305 ( .B(arr[2047]), .A(arr[2080]), .S(n2439), .Y(n412) );
  MUX2X1 U5306 ( .B(arr[1981]), .A(arr[2014]), .S(n2439), .Y(n411) );
  MUX2X1 U5307 ( .B(arr[1915]), .A(arr[1948]), .S(n2439), .Y(n415) );
  MUX2X1 U5308 ( .B(arr[1849]), .A(arr[1882]), .S(n2439), .Y(n414) );
  MUX2X1 U5309 ( .B(n413), .A(n410), .S(n2594), .Y(n424) );
  MUX2X1 U5310 ( .B(arr[1783]), .A(arr[1816]), .S(n2440), .Y(n418) );
  MUX2X1 U5311 ( .B(arr[1717]), .A(arr[1750]), .S(n2440), .Y(n417) );
  MUX2X1 U5312 ( .B(arr[1651]), .A(arr[1684]), .S(n2440), .Y(n421) );
  MUX2X1 U5313 ( .B(arr[1585]), .A(arr[1618]), .S(n2440), .Y(n420) );
  MUX2X1 U5314 ( .B(n419), .A(n416), .S(n2594), .Y(n423) );
  MUX2X1 U5315 ( .B(arr[1519]), .A(arr[1552]), .S(n2440), .Y(n427) );
  MUX2X1 U5316 ( .B(arr[1453]), .A(arr[1486]), .S(n2440), .Y(n426) );
  MUX2X1 U5317 ( .B(arr[1387]), .A(arr[1420]), .S(n2440), .Y(n430) );
  MUX2X1 U5318 ( .B(arr[1321]), .A(arr[1354]), .S(n2440), .Y(n429) );
  MUX2X1 U5319 ( .B(n428), .A(n425), .S(n2594), .Y(n439) );
  MUX2X1 U5320 ( .B(arr[1255]), .A(arr[1288]), .S(n2440), .Y(n433) );
  MUX2X1 U5321 ( .B(arr[1189]), .A(arr[1222]), .S(n2440), .Y(n432) );
  MUX2X1 U5322 ( .B(arr[1123]), .A(arr[1156]), .S(n2440), .Y(n436) );
  MUX2X1 U5323 ( .B(arr[1057]), .A(arr[1090]), .S(n2440), .Y(n435) );
  MUX2X1 U5324 ( .B(n434), .A(n431), .S(n2594), .Y(n438) );
  MUX2X1 U5325 ( .B(n437), .A(n422), .S(n2635), .Y(n471) );
  MUX2X1 U5326 ( .B(arr[991]), .A(arr[1024]), .S(n2441), .Y(n442) );
  MUX2X1 U5327 ( .B(arr[925]), .A(arr[958]), .S(n2441), .Y(n441) );
  MUX2X1 U5328 ( .B(arr[859]), .A(arr[892]), .S(n2441), .Y(n445) );
  MUX2X1 U5329 ( .B(arr[793]), .A(arr[826]), .S(n2441), .Y(n444) );
  MUX2X1 U5330 ( .B(n443), .A(n440), .S(n2595), .Y(n454) );
  MUX2X1 U5331 ( .B(arr[727]), .A(arr[760]), .S(n2441), .Y(n448) );
  MUX2X1 U5332 ( .B(arr[661]), .A(arr[694]), .S(n2441), .Y(n447) );
  MUX2X1 U5333 ( .B(arr[595]), .A(arr[628]), .S(n2441), .Y(n451) );
  MUX2X1 U5334 ( .B(arr[529]), .A(arr[562]), .S(n2441), .Y(n450) );
  MUX2X1 U5335 ( .B(n449), .A(n446), .S(n2595), .Y(n453) );
  MUX2X1 U5336 ( .B(arr[463]), .A(arr[496]), .S(n2441), .Y(n457) );
  MUX2X1 U5337 ( .B(arr[397]), .A(arr[430]), .S(n2441), .Y(n456) );
  MUX2X1 U5338 ( .B(arr[331]), .A(arr[364]), .S(n2441), .Y(n460) );
  MUX2X1 U5339 ( .B(arr[265]), .A(arr[298]), .S(n2441), .Y(n459) );
  MUX2X1 U5340 ( .B(n458), .A(n455), .S(n2595), .Y(n469) );
  MUX2X1 U5341 ( .B(arr[199]), .A(arr[232]), .S(n2442), .Y(n463) );
  MUX2X1 U5342 ( .B(arr[133]), .A(arr[166]), .S(n2442), .Y(n462) );
  MUX2X1 U5343 ( .B(arr[67]), .A(arr[100]), .S(n2442), .Y(n466) );
  MUX2X1 U5344 ( .B(arr[1]), .A(arr[34]), .S(n2442), .Y(n465) );
  MUX2X1 U5345 ( .B(n464), .A(n461), .S(n2595), .Y(n468) );
  MUX2X1 U5346 ( .B(n467), .A(n452), .S(n2635), .Y(n470) );
  MUX2X1 U5347 ( .B(arr[2048]), .A(arr[2081]), .S(n2442), .Y(n474) );
  MUX2X1 U5348 ( .B(arr[1982]), .A(arr[2015]), .S(n2442), .Y(n473) );
  MUX2X1 U5349 ( .B(arr[1916]), .A(arr[1949]), .S(n2442), .Y(n477) );
  MUX2X1 U5350 ( .B(arr[1850]), .A(arr[1883]), .S(n2442), .Y(n476) );
  MUX2X1 U5351 ( .B(n475), .A(n472), .S(n2595), .Y(n486) );
  MUX2X1 U5352 ( .B(arr[1784]), .A(arr[1817]), .S(n2442), .Y(n480) );
  MUX2X1 U5353 ( .B(arr[1718]), .A(arr[1751]), .S(n2442), .Y(n479) );
  MUX2X1 U5354 ( .B(arr[1652]), .A(arr[1685]), .S(n2442), .Y(n483) );
  MUX2X1 U5355 ( .B(arr[1586]), .A(arr[1619]), .S(n2442), .Y(n482) );
  MUX2X1 U5356 ( .B(n481), .A(n478), .S(n2595), .Y(n485) );
  MUX2X1 U5357 ( .B(arr[1520]), .A(arr[1553]), .S(n2443), .Y(n489) );
  MUX2X1 U5358 ( .B(arr[1454]), .A(arr[1487]), .S(n2443), .Y(n488) );
  MUX2X1 U5359 ( .B(arr[1388]), .A(arr[1421]), .S(n2443), .Y(n492) );
  MUX2X1 U5360 ( .B(arr[1322]), .A(arr[1355]), .S(n2443), .Y(n491) );
  MUX2X1 U5361 ( .B(n490), .A(n487), .S(n2595), .Y(n501) );
  MUX2X1 U5362 ( .B(arr[1256]), .A(arr[1289]), .S(n2443), .Y(n495) );
  MUX2X1 U5363 ( .B(arr[1190]), .A(arr[1223]), .S(n2443), .Y(n494) );
  MUX2X1 U5364 ( .B(arr[1124]), .A(arr[1157]), .S(n2443), .Y(n498) );
  MUX2X1 U5365 ( .B(arr[1058]), .A(arr[1091]), .S(n2443), .Y(n497) );
  MUX2X1 U5366 ( .B(n496), .A(n493), .S(n2595), .Y(n500) );
  MUX2X1 U5367 ( .B(n499), .A(n484), .S(n2635), .Y(n533) );
  MUX2X1 U5368 ( .B(arr[992]), .A(arr[1025]), .S(n2443), .Y(n504) );
  MUX2X1 U5369 ( .B(arr[926]), .A(arr[959]), .S(n2443), .Y(n503) );
  MUX2X1 U5370 ( .B(arr[860]), .A(arr[893]), .S(n2443), .Y(n507) );
  MUX2X1 U5371 ( .B(arr[794]), .A(arr[827]), .S(n2443), .Y(n506) );
  MUX2X1 U5372 ( .B(n505), .A(n502), .S(n2595), .Y(n516) );
  MUX2X1 U5373 ( .B(arr[728]), .A(arr[761]), .S(n2444), .Y(n510) );
  MUX2X1 U5374 ( .B(arr[662]), .A(arr[695]), .S(n2444), .Y(n509) );
  MUX2X1 U5375 ( .B(arr[596]), .A(arr[629]), .S(n2444), .Y(n513) );
  MUX2X1 U5376 ( .B(arr[530]), .A(arr[563]), .S(n2444), .Y(n512) );
  MUX2X1 U5377 ( .B(n511), .A(n508), .S(n2595), .Y(n515) );
  MUX2X1 U5378 ( .B(arr[464]), .A(arr[497]), .S(n2444), .Y(n519) );
  MUX2X1 U5379 ( .B(arr[398]), .A(arr[431]), .S(n2444), .Y(n518) );
  MUX2X1 U5380 ( .B(arr[332]), .A(arr[365]), .S(n2444), .Y(n522) );
  MUX2X1 U5381 ( .B(arr[266]), .A(arr[299]), .S(n2444), .Y(n521) );
  MUX2X1 U5382 ( .B(n520), .A(n517), .S(n2595), .Y(n531) );
  MUX2X1 U5383 ( .B(arr[200]), .A(arr[233]), .S(n2444), .Y(n525) );
  MUX2X1 U5384 ( .B(arr[134]), .A(arr[167]), .S(n2444), .Y(n524) );
  MUX2X1 U5385 ( .B(arr[68]), .A(arr[101]), .S(n2444), .Y(n528) );
  MUX2X1 U5386 ( .B(arr[2]), .A(arr[35]), .S(n2444), .Y(n527) );
  MUX2X1 U5387 ( .B(n526), .A(n523), .S(n2595), .Y(n530) );
  MUX2X1 U5388 ( .B(n529), .A(n514), .S(n2635), .Y(n532) );
  MUX2X1 U5389 ( .B(arr[2049]), .A(arr[2082]), .S(n2445), .Y(n536) );
  MUX2X1 U5390 ( .B(arr[1983]), .A(arr[2016]), .S(n2445), .Y(n535) );
  MUX2X1 U5391 ( .B(arr[1917]), .A(arr[1950]), .S(n2445), .Y(n539) );
  MUX2X1 U5392 ( .B(arr[1851]), .A(arr[1884]), .S(n2445), .Y(n538) );
  MUX2X1 U5393 ( .B(n537), .A(n534), .S(n2596), .Y(n548) );
  MUX2X1 U5394 ( .B(arr[1785]), .A(arr[1818]), .S(n2445), .Y(n542) );
  MUX2X1 U5395 ( .B(arr[1719]), .A(arr[1752]), .S(n2445), .Y(n541) );
  MUX2X1 U5396 ( .B(arr[1653]), .A(arr[1686]), .S(n2445), .Y(n545) );
  MUX2X1 U5397 ( .B(arr[1587]), .A(arr[1620]), .S(n2445), .Y(n544) );
  MUX2X1 U5398 ( .B(n543), .A(n540), .S(n2596), .Y(n547) );
  MUX2X1 U5399 ( .B(arr[1521]), .A(arr[1554]), .S(n2445), .Y(n551) );
  MUX2X1 U5400 ( .B(arr[1455]), .A(arr[1488]), .S(n2445), .Y(n550) );
  MUX2X1 U5401 ( .B(arr[1389]), .A(arr[1422]), .S(n2445), .Y(n554) );
  MUX2X1 U5402 ( .B(arr[1323]), .A(arr[1356]), .S(n2445), .Y(n553) );
  MUX2X1 U5403 ( .B(n552), .A(n549), .S(n2596), .Y(n563) );
  MUX2X1 U5404 ( .B(arr[1257]), .A(arr[1290]), .S(n2446), .Y(n557) );
  MUX2X1 U5405 ( .B(arr[1191]), .A(arr[1224]), .S(n2446), .Y(n556) );
  MUX2X1 U5406 ( .B(arr[1125]), .A(arr[1158]), .S(n2446), .Y(n560) );
  MUX2X1 U5407 ( .B(arr[1059]), .A(arr[1092]), .S(n2446), .Y(n559) );
  MUX2X1 U5408 ( .B(n558), .A(n555), .S(n2596), .Y(n562) );
  MUX2X1 U5409 ( .B(n561), .A(n546), .S(n2636), .Y(n595) );
  MUX2X1 U5410 ( .B(arr[993]), .A(arr[1026]), .S(n2446), .Y(n566) );
  MUX2X1 U5411 ( .B(arr[927]), .A(arr[960]), .S(n2446), .Y(n565) );
  MUX2X1 U5412 ( .B(arr[861]), .A(arr[894]), .S(n2446), .Y(n569) );
  MUX2X1 U5413 ( .B(arr[795]), .A(arr[828]), .S(n2446), .Y(n568) );
  MUX2X1 U5414 ( .B(n567), .A(n564), .S(n2596), .Y(n578) );
  MUX2X1 U5415 ( .B(arr[729]), .A(arr[762]), .S(n2446), .Y(n572) );
  MUX2X1 U5416 ( .B(arr[663]), .A(arr[696]), .S(n2446), .Y(n571) );
  MUX2X1 U5417 ( .B(arr[597]), .A(arr[630]), .S(n2446), .Y(n575) );
  MUX2X1 U5418 ( .B(arr[531]), .A(arr[564]), .S(n2446), .Y(n574) );
  MUX2X1 U5419 ( .B(n573), .A(n570), .S(n2596), .Y(n577) );
  MUX2X1 U5420 ( .B(arr[465]), .A(arr[498]), .S(n2447), .Y(n581) );
  MUX2X1 U5421 ( .B(arr[399]), .A(arr[432]), .S(n2447), .Y(n580) );
  MUX2X1 U5422 ( .B(arr[333]), .A(arr[366]), .S(n2447), .Y(n584) );
  MUX2X1 U5423 ( .B(arr[267]), .A(arr[300]), .S(n2447), .Y(n583) );
  MUX2X1 U5424 ( .B(n582), .A(n579), .S(n2596), .Y(n593) );
  MUX2X1 U5425 ( .B(arr[201]), .A(arr[234]), .S(n2447), .Y(n587) );
  MUX2X1 U5426 ( .B(arr[135]), .A(arr[168]), .S(n2447), .Y(n586) );
  MUX2X1 U5427 ( .B(arr[69]), .A(arr[102]), .S(n2447), .Y(n590) );
  MUX2X1 U5428 ( .B(arr[3]), .A(arr[36]), .S(n2447), .Y(n589) );
  MUX2X1 U5429 ( .B(n588), .A(n585), .S(n2596), .Y(n592) );
  MUX2X1 U5430 ( .B(n591), .A(n576), .S(n2636), .Y(n594) );
  MUX2X1 U5431 ( .B(arr[2050]), .A(arr[2083]), .S(n2447), .Y(n598) );
  MUX2X1 U5432 ( .B(arr[1984]), .A(arr[2017]), .S(n2447), .Y(n597) );
  MUX2X1 U5433 ( .B(arr[1918]), .A(arr[1951]), .S(n2447), .Y(n601) );
  MUX2X1 U5434 ( .B(arr[1852]), .A(arr[1885]), .S(n2447), .Y(n600) );
  MUX2X1 U5435 ( .B(n599), .A(n596), .S(n2596), .Y(n610) );
  MUX2X1 U5436 ( .B(arr[1786]), .A(arr[1819]), .S(n2448), .Y(n604) );
  MUX2X1 U5437 ( .B(arr[1720]), .A(arr[1753]), .S(n2448), .Y(n603) );
  MUX2X1 U5438 ( .B(arr[1654]), .A(arr[1687]), .S(n2448), .Y(n607) );
  MUX2X1 U5439 ( .B(arr[1588]), .A(arr[1621]), .S(n2448), .Y(n606) );
  MUX2X1 U5440 ( .B(n605), .A(n602), .S(n2596), .Y(n609) );
  MUX2X1 U5441 ( .B(arr[1522]), .A(arr[1555]), .S(n2448), .Y(n613) );
  MUX2X1 U5442 ( .B(arr[1456]), .A(arr[1489]), .S(n2448), .Y(n612) );
  MUX2X1 U5443 ( .B(arr[1390]), .A(arr[1423]), .S(n2448), .Y(n616) );
  MUX2X1 U5444 ( .B(arr[1324]), .A(arr[1357]), .S(n2448), .Y(n615) );
  MUX2X1 U5445 ( .B(n614), .A(n611), .S(n2596), .Y(n625) );
  MUX2X1 U5446 ( .B(arr[1258]), .A(arr[1291]), .S(n2448), .Y(n619) );
  MUX2X1 U5447 ( .B(arr[1192]), .A(arr[1225]), .S(n2448), .Y(n618) );
  MUX2X1 U5448 ( .B(arr[1126]), .A(arr[1159]), .S(n2448), .Y(n622) );
  MUX2X1 U5449 ( .B(arr[1060]), .A(arr[1093]), .S(n2448), .Y(n621) );
  MUX2X1 U5450 ( .B(n620), .A(n617), .S(n2596), .Y(n624) );
  MUX2X1 U5451 ( .B(n623), .A(n608), .S(n2636), .Y(n657) );
  MUX2X1 U5452 ( .B(arr[994]), .A(arr[1027]), .S(n2449), .Y(n628) );
  MUX2X1 U5453 ( .B(arr[928]), .A(arr[961]), .S(n2449), .Y(n627) );
  MUX2X1 U5454 ( .B(arr[862]), .A(arr[895]), .S(n2449), .Y(n631) );
  MUX2X1 U5455 ( .B(arr[796]), .A(arr[829]), .S(n2449), .Y(n630) );
  MUX2X1 U5456 ( .B(n629), .A(n626), .S(n2597), .Y(n640) );
  MUX2X1 U5457 ( .B(arr[730]), .A(arr[763]), .S(n2449), .Y(n634) );
  MUX2X1 U5458 ( .B(arr[664]), .A(arr[697]), .S(n2449), .Y(n633) );
  MUX2X1 U5459 ( .B(arr[598]), .A(arr[631]), .S(n2449), .Y(n637) );
  MUX2X1 U5460 ( .B(arr[532]), .A(arr[565]), .S(n2449), .Y(n636) );
  MUX2X1 U5461 ( .B(n635), .A(n632), .S(n2597), .Y(n639) );
  MUX2X1 U5462 ( .B(arr[466]), .A(arr[499]), .S(n2449), .Y(n643) );
  MUX2X1 U5463 ( .B(arr[400]), .A(arr[433]), .S(n2449), .Y(n642) );
  MUX2X1 U5464 ( .B(arr[334]), .A(arr[367]), .S(n2449), .Y(n646) );
  MUX2X1 U5465 ( .B(arr[268]), .A(arr[301]), .S(n2449), .Y(n645) );
  MUX2X1 U5466 ( .B(n644), .A(n641), .S(n2597), .Y(n655) );
  MUX2X1 U5467 ( .B(arr[202]), .A(arr[235]), .S(n2450), .Y(n649) );
  MUX2X1 U5468 ( .B(arr[136]), .A(arr[169]), .S(n2450), .Y(n648) );
  MUX2X1 U5469 ( .B(arr[70]), .A(arr[103]), .S(n2450), .Y(n652) );
  MUX2X1 U5470 ( .B(arr[4]), .A(arr[37]), .S(n2450), .Y(n651) );
  MUX2X1 U5471 ( .B(n650), .A(n647), .S(n2597), .Y(n654) );
  MUX2X1 U5472 ( .B(n653), .A(n638), .S(n2636), .Y(n656) );
  MUX2X1 U5473 ( .B(arr[2051]), .A(arr[2084]), .S(n2450), .Y(n660) );
  MUX2X1 U5474 ( .B(arr[1985]), .A(arr[2018]), .S(n2450), .Y(n659) );
  MUX2X1 U5475 ( .B(arr[1919]), .A(arr[1952]), .S(n2450), .Y(n663) );
  MUX2X1 U5476 ( .B(arr[1853]), .A(arr[1886]), .S(n2450), .Y(n662) );
  MUX2X1 U5477 ( .B(n661), .A(n658), .S(n2597), .Y(n672) );
  MUX2X1 U5478 ( .B(arr[1787]), .A(arr[1820]), .S(n2450), .Y(n666) );
  MUX2X1 U5479 ( .B(arr[1721]), .A(arr[1754]), .S(n2450), .Y(n665) );
  MUX2X1 U5480 ( .B(arr[1655]), .A(arr[1688]), .S(n2450), .Y(n669) );
  MUX2X1 U5481 ( .B(arr[1589]), .A(arr[1622]), .S(n2450), .Y(n668) );
  MUX2X1 U5482 ( .B(n667), .A(n664), .S(n2597), .Y(n671) );
  MUX2X1 U5483 ( .B(arr[1523]), .A(arr[1556]), .S(n2451), .Y(n675) );
  MUX2X1 U5484 ( .B(arr[1457]), .A(arr[1490]), .S(n2451), .Y(n674) );
  MUX2X1 U5485 ( .B(arr[1391]), .A(arr[1424]), .S(n2451), .Y(n678) );
  MUX2X1 U5486 ( .B(arr[1325]), .A(arr[1358]), .S(n2451), .Y(n677) );
  MUX2X1 U5487 ( .B(n676), .A(n673), .S(n2597), .Y(n687) );
  MUX2X1 U5488 ( .B(arr[1259]), .A(arr[1292]), .S(n2451), .Y(n681) );
  MUX2X1 U5489 ( .B(arr[1193]), .A(arr[1226]), .S(n2451), .Y(n680) );
  MUX2X1 U5490 ( .B(arr[1127]), .A(arr[1160]), .S(n2451), .Y(n684) );
  MUX2X1 U5491 ( .B(arr[1061]), .A(arr[1094]), .S(n2451), .Y(n683) );
  MUX2X1 U5492 ( .B(n682), .A(n679), .S(n2597), .Y(n686) );
  MUX2X1 U5493 ( .B(n685), .A(n670), .S(n2636), .Y(n719) );
  MUX2X1 U5494 ( .B(arr[995]), .A(arr[1028]), .S(n2451), .Y(n690) );
  MUX2X1 U5495 ( .B(arr[929]), .A(arr[962]), .S(n2451), .Y(n689) );
  MUX2X1 U5496 ( .B(arr[863]), .A(arr[896]), .S(n2451), .Y(n693) );
  MUX2X1 U5497 ( .B(arr[797]), .A(arr[830]), .S(n2451), .Y(n692) );
  MUX2X1 U5498 ( .B(n691), .A(n688), .S(n2597), .Y(n702) );
  MUX2X1 U5499 ( .B(arr[731]), .A(arr[764]), .S(n2452), .Y(n696) );
  MUX2X1 U5500 ( .B(arr[665]), .A(arr[698]), .S(n2452), .Y(n695) );
  MUX2X1 U5501 ( .B(arr[599]), .A(arr[632]), .S(n2452), .Y(n699) );
  MUX2X1 U5502 ( .B(arr[533]), .A(arr[566]), .S(n2452), .Y(n698) );
  MUX2X1 U5503 ( .B(n697), .A(n694), .S(n2597), .Y(n701) );
  MUX2X1 U5504 ( .B(arr[467]), .A(arr[500]), .S(n2452), .Y(n705) );
  MUX2X1 U5505 ( .B(arr[401]), .A(arr[434]), .S(n2452), .Y(n704) );
  MUX2X1 U5506 ( .B(arr[335]), .A(arr[368]), .S(n2452), .Y(n708) );
  MUX2X1 U5507 ( .B(arr[269]), .A(arr[302]), .S(n2452), .Y(n707) );
  MUX2X1 U5508 ( .B(n706), .A(n703), .S(n2597), .Y(n717) );
  MUX2X1 U5509 ( .B(arr[203]), .A(arr[236]), .S(n2452), .Y(n711) );
  MUX2X1 U5510 ( .B(arr[137]), .A(arr[170]), .S(n2452), .Y(n710) );
  MUX2X1 U5511 ( .B(arr[71]), .A(arr[104]), .S(n2452), .Y(n714) );
  MUX2X1 U5512 ( .B(arr[5]), .A(arr[38]), .S(n2452), .Y(n713) );
  MUX2X1 U5513 ( .B(n712), .A(n709), .S(n2597), .Y(n716) );
  MUX2X1 U5514 ( .B(n715), .A(n700), .S(n2636), .Y(n718) );
  MUX2X1 U5515 ( .B(arr[2052]), .A(arr[2085]), .S(n2453), .Y(n722) );
  MUX2X1 U5516 ( .B(arr[1986]), .A(arr[2019]), .S(n2453), .Y(n721) );
  MUX2X1 U5517 ( .B(arr[1920]), .A(arr[1953]), .S(n2453), .Y(n725) );
  MUX2X1 U5518 ( .B(arr[1854]), .A(arr[1887]), .S(n2453), .Y(n724) );
  MUX2X1 U5519 ( .B(n723), .A(n720), .S(n2598), .Y(n734) );
  MUX2X1 U5520 ( .B(arr[1788]), .A(arr[1821]), .S(n2453), .Y(n728) );
  MUX2X1 U5521 ( .B(arr[1722]), .A(arr[1755]), .S(n2453), .Y(n727) );
  MUX2X1 U5522 ( .B(arr[1656]), .A(arr[1689]), .S(n2453), .Y(n731) );
  MUX2X1 U5523 ( .B(arr[1590]), .A(arr[1623]), .S(n2453), .Y(n730) );
  MUX2X1 U5524 ( .B(n729), .A(n726), .S(n2598), .Y(n733) );
  MUX2X1 U5525 ( .B(arr[1524]), .A(arr[1557]), .S(n2453), .Y(n737) );
  MUX2X1 U5526 ( .B(arr[1458]), .A(arr[1491]), .S(n2453), .Y(n736) );
  MUX2X1 U5527 ( .B(arr[1392]), .A(arr[1425]), .S(n2453), .Y(n740) );
  MUX2X1 U5528 ( .B(arr[1326]), .A(arr[1359]), .S(n2453), .Y(n739) );
  MUX2X1 U5529 ( .B(n738), .A(n735), .S(n2598), .Y(n749) );
  MUX2X1 U5530 ( .B(arr[1260]), .A(arr[1293]), .S(n2454), .Y(n743) );
  MUX2X1 U5531 ( .B(arr[1194]), .A(arr[1227]), .S(n2454), .Y(n742) );
  MUX2X1 U5532 ( .B(arr[1128]), .A(arr[1161]), .S(n2454), .Y(n746) );
  MUX2X1 U5533 ( .B(arr[1062]), .A(arr[1095]), .S(n2454), .Y(n745) );
  MUX2X1 U5534 ( .B(n744), .A(n741), .S(n2598), .Y(n748) );
  MUX2X1 U5535 ( .B(n747), .A(n732), .S(n2636), .Y(n781) );
  MUX2X1 U5536 ( .B(arr[996]), .A(arr[1029]), .S(n2454), .Y(n752) );
  MUX2X1 U5537 ( .B(arr[930]), .A(arr[963]), .S(n2454), .Y(n751) );
  MUX2X1 U5538 ( .B(arr[864]), .A(arr[897]), .S(n2454), .Y(n755) );
  MUX2X1 U5539 ( .B(arr[798]), .A(arr[831]), .S(n2454), .Y(n754) );
  MUX2X1 U5540 ( .B(n753), .A(n750), .S(n2598), .Y(n764) );
  MUX2X1 U5541 ( .B(arr[732]), .A(arr[765]), .S(n2454), .Y(n758) );
  MUX2X1 U5542 ( .B(arr[666]), .A(arr[699]), .S(n2454), .Y(n757) );
  MUX2X1 U5543 ( .B(arr[600]), .A(arr[633]), .S(n2454), .Y(n761) );
  MUX2X1 U5544 ( .B(arr[534]), .A(arr[567]), .S(n2454), .Y(n760) );
  MUX2X1 U5545 ( .B(n759), .A(n756), .S(n2598), .Y(n763) );
  MUX2X1 U5546 ( .B(arr[468]), .A(arr[501]), .S(n2455), .Y(n767) );
  MUX2X1 U5547 ( .B(arr[402]), .A(arr[435]), .S(n2455), .Y(n766) );
  MUX2X1 U5548 ( .B(arr[336]), .A(arr[369]), .S(n2455), .Y(n770) );
  MUX2X1 U5549 ( .B(arr[270]), .A(arr[303]), .S(n2455), .Y(n769) );
  MUX2X1 U5550 ( .B(n768), .A(n765), .S(n2598), .Y(n779) );
  MUX2X1 U5551 ( .B(arr[204]), .A(arr[237]), .S(n2455), .Y(n773) );
  MUX2X1 U5552 ( .B(arr[138]), .A(arr[171]), .S(n2455), .Y(n772) );
  MUX2X1 U5553 ( .B(arr[72]), .A(arr[105]), .S(n2455), .Y(n776) );
  MUX2X1 U5554 ( .B(arr[6]), .A(arr[39]), .S(n2455), .Y(n775) );
  MUX2X1 U5555 ( .B(n774), .A(n771), .S(n2598), .Y(n778) );
  MUX2X1 U5556 ( .B(n777), .A(n762), .S(n2636), .Y(n780) );
  MUX2X1 U5557 ( .B(arr[2053]), .A(arr[2086]), .S(n2455), .Y(n784) );
  MUX2X1 U5558 ( .B(arr[1987]), .A(arr[2020]), .S(n2455), .Y(n783) );
  MUX2X1 U5559 ( .B(arr[1921]), .A(arr[1954]), .S(n2455), .Y(n787) );
  MUX2X1 U5560 ( .B(arr[1855]), .A(arr[1888]), .S(n2455), .Y(n786) );
  MUX2X1 U5561 ( .B(n785), .A(n782), .S(n2598), .Y(n796) );
  MUX2X1 U5562 ( .B(arr[1789]), .A(arr[1822]), .S(n2456), .Y(n790) );
  MUX2X1 U5563 ( .B(arr[1723]), .A(arr[1756]), .S(n2456), .Y(n789) );
  MUX2X1 U5564 ( .B(arr[1657]), .A(arr[1690]), .S(n2456), .Y(n793) );
  MUX2X1 U5565 ( .B(arr[1591]), .A(arr[1624]), .S(n2456), .Y(n792) );
  MUX2X1 U5566 ( .B(n791), .A(n788), .S(n2598), .Y(n795) );
  MUX2X1 U5567 ( .B(arr[1525]), .A(arr[1558]), .S(n2456), .Y(n799) );
  MUX2X1 U5568 ( .B(arr[1459]), .A(arr[1492]), .S(n2456), .Y(n798) );
  MUX2X1 U5569 ( .B(arr[1393]), .A(arr[1426]), .S(n2456), .Y(n802) );
  MUX2X1 U5570 ( .B(arr[1327]), .A(arr[1360]), .S(n2456), .Y(n801) );
  MUX2X1 U5571 ( .B(n800), .A(n797), .S(n2598), .Y(n811) );
  MUX2X1 U5572 ( .B(arr[1261]), .A(arr[1294]), .S(n2456), .Y(n805) );
  MUX2X1 U5573 ( .B(arr[1195]), .A(arr[1228]), .S(n2456), .Y(n804) );
  MUX2X1 U5574 ( .B(arr[1129]), .A(arr[1162]), .S(n2456), .Y(n808) );
  MUX2X1 U5575 ( .B(arr[1063]), .A(arr[1096]), .S(n2456), .Y(n807) );
  MUX2X1 U5576 ( .B(n806), .A(n803), .S(n2598), .Y(n810) );
  MUX2X1 U5577 ( .B(n809), .A(n794), .S(n2636), .Y(n843) );
  MUX2X1 U5578 ( .B(arr[997]), .A(arr[1030]), .S(n2457), .Y(n814) );
  MUX2X1 U5579 ( .B(arr[931]), .A(arr[964]), .S(n2457), .Y(n813) );
  MUX2X1 U5580 ( .B(arr[865]), .A(arr[898]), .S(n2457), .Y(n817) );
  MUX2X1 U5581 ( .B(arr[799]), .A(arr[832]), .S(n2457), .Y(n816) );
  MUX2X1 U5582 ( .B(n815), .A(n812), .S(n2599), .Y(n826) );
  MUX2X1 U5583 ( .B(arr[733]), .A(arr[766]), .S(n2457), .Y(n820) );
  MUX2X1 U5584 ( .B(arr[667]), .A(arr[700]), .S(n2457), .Y(n819) );
  MUX2X1 U5585 ( .B(arr[601]), .A(arr[634]), .S(n2457), .Y(n823) );
  MUX2X1 U5586 ( .B(arr[535]), .A(arr[568]), .S(n2457), .Y(n822) );
  MUX2X1 U5587 ( .B(n821), .A(n818), .S(n2599), .Y(n825) );
  MUX2X1 U5588 ( .B(arr[469]), .A(arr[502]), .S(n2457), .Y(n829) );
  MUX2X1 U5589 ( .B(arr[403]), .A(arr[436]), .S(n2457), .Y(n828) );
  MUX2X1 U5590 ( .B(arr[337]), .A(arr[370]), .S(n2457), .Y(n832) );
  MUX2X1 U5591 ( .B(arr[271]), .A(arr[304]), .S(n2457), .Y(n831) );
  MUX2X1 U5592 ( .B(n830), .A(n827), .S(n2599), .Y(n841) );
  MUX2X1 U5593 ( .B(arr[205]), .A(arr[238]), .S(n2458), .Y(n835) );
  MUX2X1 U5594 ( .B(arr[139]), .A(arr[172]), .S(n2458), .Y(n834) );
  MUX2X1 U5595 ( .B(arr[73]), .A(arr[106]), .S(n2458), .Y(n838) );
  MUX2X1 U5596 ( .B(arr[7]), .A(arr[40]), .S(n2458), .Y(n837) );
  MUX2X1 U5597 ( .B(n836), .A(n833), .S(n2599), .Y(n840) );
  MUX2X1 U5598 ( .B(n839), .A(n824), .S(n2636), .Y(n842) );
  MUX2X1 U5599 ( .B(arr[2054]), .A(arr[2087]), .S(n2458), .Y(n846) );
  MUX2X1 U5600 ( .B(arr[1988]), .A(arr[2021]), .S(n2458), .Y(n845) );
  MUX2X1 U5601 ( .B(arr[1922]), .A(arr[1955]), .S(n2458), .Y(n849) );
  MUX2X1 U5602 ( .B(arr[1856]), .A(arr[1889]), .S(n2458), .Y(n848) );
  MUX2X1 U5603 ( .B(n847), .A(n844), .S(n2599), .Y(n858) );
  MUX2X1 U5604 ( .B(arr[1790]), .A(arr[1823]), .S(n2458), .Y(n852) );
  MUX2X1 U5605 ( .B(arr[1724]), .A(arr[1757]), .S(n2458), .Y(n851) );
  MUX2X1 U5606 ( .B(arr[1658]), .A(arr[1691]), .S(n2458), .Y(n855) );
  MUX2X1 U5607 ( .B(arr[1592]), .A(arr[1625]), .S(n2458), .Y(n854) );
  MUX2X1 U5608 ( .B(n853), .A(n850), .S(n2599), .Y(n857) );
  MUX2X1 U5609 ( .B(arr[1526]), .A(arr[1559]), .S(n2459), .Y(n861) );
  MUX2X1 U5610 ( .B(arr[1460]), .A(arr[1493]), .S(n2459), .Y(n860) );
  MUX2X1 U5611 ( .B(arr[1394]), .A(arr[1427]), .S(n2459), .Y(n864) );
  MUX2X1 U5612 ( .B(arr[1328]), .A(arr[1361]), .S(n2459), .Y(n863) );
  MUX2X1 U5613 ( .B(n862), .A(n859), .S(n2599), .Y(n873) );
  MUX2X1 U5614 ( .B(arr[1262]), .A(arr[1295]), .S(n2459), .Y(n867) );
  MUX2X1 U5615 ( .B(arr[1196]), .A(arr[1229]), .S(n2459), .Y(n866) );
  MUX2X1 U5616 ( .B(arr[1130]), .A(arr[1163]), .S(n2459), .Y(n870) );
  MUX2X1 U5617 ( .B(arr[1064]), .A(arr[1097]), .S(n2459), .Y(n869) );
  MUX2X1 U5618 ( .B(n868), .A(n865), .S(n2599), .Y(n872) );
  MUX2X1 U5619 ( .B(n871), .A(n856), .S(n2636), .Y(n905) );
  MUX2X1 U5620 ( .B(arr[998]), .A(arr[1031]), .S(n2459), .Y(n876) );
  MUX2X1 U5621 ( .B(arr[932]), .A(arr[965]), .S(n2459), .Y(n875) );
  MUX2X1 U5622 ( .B(arr[866]), .A(arr[899]), .S(n2459), .Y(n879) );
  MUX2X1 U5623 ( .B(arr[800]), .A(arr[833]), .S(n2459), .Y(n878) );
  MUX2X1 U5624 ( .B(n877), .A(n874), .S(n2599), .Y(n888) );
  MUX2X1 U5625 ( .B(arr[734]), .A(arr[767]), .S(n2460), .Y(n882) );
  MUX2X1 U5626 ( .B(arr[668]), .A(arr[701]), .S(n2460), .Y(n881) );
  MUX2X1 U5627 ( .B(arr[602]), .A(arr[635]), .S(n2460), .Y(n885) );
  MUX2X1 U5628 ( .B(arr[536]), .A(arr[569]), .S(n2460), .Y(n884) );
  MUX2X1 U5629 ( .B(n883), .A(n880), .S(n2599), .Y(n887) );
  MUX2X1 U5630 ( .B(arr[470]), .A(arr[503]), .S(n2460), .Y(n891) );
  MUX2X1 U5631 ( .B(arr[404]), .A(arr[437]), .S(n2460), .Y(n890) );
  MUX2X1 U5632 ( .B(arr[338]), .A(arr[371]), .S(n2460), .Y(n894) );
  MUX2X1 U5633 ( .B(arr[272]), .A(arr[305]), .S(n2460), .Y(n893) );
  MUX2X1 U5634 ( .B(n892), .A(n889), .S(n2599), .Y(n903) );
  MUX2X1 U5635 ( .B(arr[206]), .A(arr[239]), .S(n2460), .Y(n897) );
  MUX2X1 U5636 ( .B(arr[140]), .A(arr[173]), .S(n2460), .Y(n896) );
  MUX2X1 U5637 ( .B(arr[74]), .A(arr[107]), .S(n2460), .Y(n900) );
  MUX2X1 U5638 ( .B(arr[8]), .A(arr[41]), .S(n2460), .Y(n899) );
  MUX2X1 U5639 ( .B(n898), .A(n895), .S(n2599), .Y(n902) );
  MUX2X1 U5640 ( .B(n901), .A(n886), .S(n2636), .Y(n904) );
  MUX2X1 U5641 ( .B(arr[2055]), .A(arr[2088]), .S(n2461), .Y(n908) );
  MUX2X1 U5642 ( .B(arr[1989]), .A(arr[2022]), .S(n2461), .Y(n907) );
  MUX2X1 U5643 ( .B(arr[1923]), .A(arr[1956]), .S(n2461), .Y(n911) );
  MUX2X1 U5644 ( .B(arr[1857]), .A(arr[1890]), .S(n2461), .Y(n910) );
  MUX2X1 U5645 ( .B(n909), .A(n906), .S(n2600), .Y(n920) );
  MUX2X1 U5646 ( .B(arr[1791]), .A(arr[1824]), .S(n2461), .Y(n914) );
  MUX2X1 U5647 ( .B(arr[1725]), .A(arr[1758]), .S(n2461), .Y(n913) );
  MUX2X1 U5648 ( .B(arr[1659]), .A(arr[1692]), .S(n2461), .Y(n917) );
  MUX2X1 U5649 ( .B(arr[1593]), .A(arr[1626]), .S(n2461), .Y(n916) );
  MUX2X1 U5650 ( .B(n915), .A(n912), .S(n2600), .Y(n919) );
  MUX2X1 U5651 ( .B(arr[1527]), .A(arr[1560]), .S(n2461), .Y(n923) );
  MUX2X1 U5652 ( .B(arr[1461]), .A(arr[1494]), .S(n2461), .Y(n922) );
  MUX2X1 U5653 ( .B(arr[1395]), .A(arr[1428]), .S(n2461), .Y(n926) );
  MUX2X1 U5654 ( .B(arr[1329]), .A(arr[1362]), .S(n2461), .Y(n925) );
  MUX2X1 U5655 ( .B(n924), .A(n921), .S(n2600), .Y(n935) );
  MUX2X1 U5656 ( .B(arr[1263]), .A(arr[1296]), .S(n2462), .Y(n929) );
  MUX2X1 U5657 ( .B(arr[1197]), .A(arr[1230]), .S(n2462), .Y(n928) );
  MUX2X1 U5658 ( .B(arr[1131]), .A(arr[1164]), .S(n2462), .Y(n932) );
  MUX2X1 U5659 ( .B(arr[1065]), .A(arr[1098]), .S(n2462), .Y(n931) );
  MUX2X1 U5660 ( .B(n930), .A(n927), .S(n2600), .Y(n934) );
  MUX2X1 U5661 ( .B(n933), .A(n918), .S(n2637), .Y(n967) );
  MUX2X1 U5662 ( .B(arr[999]), .A(arr[1032]), .S(n2462), .Y(n938) );
  MUX2X1 U5663 ( .B(arr[933]), .A(arr[966]), .S(n2462), .Y(n937) );
  MUX2X1 U5664 ( .B(arr[867]), .A(arr[900]), .S(n2462), .Y(n941) );
  MUX2X1 U5665 ( .B(arr[801]), .A(arr[834]), .S(n2462), .Y(n940) );
  MUX2X1 U5666 ( .B(n939), .A(n936), .S(n2600), .Y(n950) );
  MUX2X1 U5667 ( .B(arr[735]), .A(arr[768]), .S(n2462), .Y(n944) );
  MUX2X1 U5668 ( .B(arr[669]), .A(arr[702]), .S(n2462), .Y(n943) );
  MUX2X1 U5669 ( .B(arr[603]), .A(arr[636]), .S(n2462), .Y(n947) );
  MUX2X1 U5670 ( .B(arr[537]), .A(arr[570]), .S(n2462), .Y(n946) );
  MUX2X1 U5671 ( .B(n945), .A(n942), .S(n2600), .Y(n949) );
  MUX2X1 U5672 ( .B(arr[471]), .A(arr[504]), .S(n2463), .Y(n953) );
  MUX2X1 U5673 ( .B(arr[405]), .A(arr[438]), .S(n2463), .Y(n952) );
  MUX2X1 U5674 ( .B(arr[339]), .A(arr[372]), .S(n2463), .Y(n956) );
  MUX2X1 U5675 ( .B(arr[273]), .A(arr[306]), .S(n2463), .Y(n955) );
  MUX2X1 U5676 ( .B(n954), .A(n951), .S(n2600), .Y(n965) );
  MUX2X1 U5677 ( .B(arr[207]), .A(arr[240]), .S(n2463), .Y(n959) );
  MUX2X1 U5678 ( .B(arr[141]), .A(arr[174]), .S(n2463), .Y(n958) );
  MUX2X1 U5679 ( .B(arr[75]), .A(arr[108]), .S(n2463), .Y(n962) );
  MUX2X1 U5680 ( .B(arr[9]), .A(arr[42]), .S(n2463), .Y(n961) );
  MUX2X1 U5681 ( .B(n960), .A(n957), .S(n2600), .Y(n964) );
  MUX2X1 U5682 ( .B(n963), .A(n948), .S(n2637), .Y(n966) );
  MUX2X1 U5683 ( .B(arr[2056]), .A(arr[2089]), .S(n2463), .Y(n970) );
  MUX2X1 U5684 ( .B(arr[1990]), .A(arr[2023]), .S(n2463), .Y(n969) );
  MUX2X1 U5685 ( .B(arr[1924]), .A(arr[1957]), .S(n2463), .Y(n973) );
  MUX2X1 U5686 ( .B(arr[1858]), .A(arr[1891]), .S(n2463), .Y(n972) );
  MUX2X1 U5687 ( .B(n971), .A(n968), .S(n2600), .Y(n982) );
  MUX2X1 U5688 ( .B(arr[1792]), .A(arr[1825]), .S(n2464), .Y(n976) );
  MUX2X1 U5689 ( .B(arr[1726]), .A(arr[1759]), .S(n2464), .Y(n975) );
  MUX2X1 U5690 ( .B(arr[1660]), .A(arr[1693]), .S(n2464), .Y(n979) );
  MUX2X1 U5691 ( .B(arr[1594]), .A(arr[1627]), .S(n2464), .Y(n978) );
  MUX2X1 U5692 ( .B(n977), .A(n974), .S(n2600), .Y(n981) );
  MUX2X1 U5693 ( .B(arr[1528]), .A(arr[1561]), .S(n2464), .Y(n985) );
  MUX2X1 U5694 ( .B(arr[1462]), .A(arr[1495]), .S(n2464), .Y(n984) );
  MUX2X1 U5695 ( .B(arr[1396]), .A(arr[1429]), .S(n2464), .Y(n988) );
  MUX2X1 U5696 ( .B(arr[1330]), .A(arr[1363]), .S(n2464), .Y(n987) );
  MUX2X1 U5697 ( .B(n986), .A(n983), .S(n2600), .Y(n997) );
  MUX2X1 U5698 ( .B(arr[1264]), .A(arr[1297]), .S(n2464), .Y(n991) );
  MUX2X1 U5699 ( .B(arr[1198]), .A(arr[1231]), .S(n2464), .Y(n990) );
  MUX2X1 U5700 ( .B(arr[1132]), .A(arr[1165]), .S(n2464), .Y(n994) );
  MUX2X1 U5701 ( .B(arr[1066]), .A(arr[1099]), .S(n2464), .Y(n993) );
  MUX2X1 U5702 ( .B(n992), .A(n989), .S(n2600), .Y(n996) );
  MUX2X1 U5703 ( .B(n995), .A(n980), .S(n2637), .Y(n1029) );
  MUX2X1 U5704 ( .B(arr[1000]), .A(arr[1033]), .S(n2465), .Y(n1000) );
  MUX2X1 U5705 ( .B(arr[934]), .A(arr[967]), .S(n2465), .Y(n999) );
  MUX2X1 U5706 ( .B(arr[868]), .A(arr[901]), .S(n2465), .Y(n1003) );
  MUX2X1 U5707 ( .B(arr[802]), .A(arr[835]), .S(n2465), .Y(n1002) );
  MUX2X1 U5708 ( .B(n1001), .A(n998), .S(n2601), .Y(n1012) );
  MUX2X1 U5709 ( .B(arr[736]), .A(arr[769]), .S(n2465), .Y(n1006) );
  MUX2X1 U5710 ( .B(arr[670]), .A(arr[703]), .S(n2465), .Y(n1005) );
  MUX2X1 U5711 ( .B(arr[604]), .A(arr[637]), .S(n2465), .Y(n1009) );
  MUX2X1 U5712 ( .B(arr[538]), .A(arr[571]), .S(n2465), .Y(n1008) );
  MUX2X1 U5713 ( .B(n1007), .A(n1004), .S(n2601), .Y(n1011) );
  MUX2X1 U5714 ( .B(arr[472]), .A(arr[505]), .S(n2465), .Y(n1015) );
  MUX2X1 U5715 ( .B(arr[406]), .A(arr[439]), .S(n2465), .Y(n1014) );
  MUX2X1 U5716 ( .B(arr[340]), .A(arr[373]), .S(n2465), .Y(n1018) );
  MUX2X1 U5717 ( .B(arr[274]), .A(arr[307]), .S(n2465), .Y(n1017) );
  MUX2X1 U5718 ( .B(n1016), .A(n1013), .S(n2601), .Y(n1027) );
  MUX2X1 U5719 ( .B(arr[208]), .A(arr[241]), .S(n2466), .Y(n1021) );
  MUX2X1 U5720 ( .B(arr[142]), .A(arr[175]), .S(n2466), .Y(n1020) );
  MUX2X1 U5721 ( .B(arr[76]), .A(arr[109]), .S(n2466), .Y(n1024) );
  MUX2X1 U5722 ( .B(arr[10]), .A(arr[43]), .S(n2466), .Y(n1023) );
  MUX2X1 U5723 ( .B(n1022), .A(n1019), .S(n2601), .Y(n1026) );
  MUX2X1 U5724 ( .B(n1025), .A(n1010), .S(n2637), .Y(n1028) );
  MUX2X1 U5725 ( .B(arr[2057]), .A(arr[2090]), .S(n2466), .Y(n1032) );
  MUX2X1 U5726 ( .B(arr[1991]), .A(arr[2024]), .S(n2466), .Y(n1031) );
  MUX2X1 U5727 ( .B(arr[1925]), .A(arr[1958]), .S(n2466), .Y(n1035) );
  MUX2X1 U5728 ( .B(arr[1859]), .A(arr[1892]), .S(n2466), .Y(n1034) );
  MUX2X1 U5729 ( .B(n1033), .A(n1030), .S(n2601), .Y(n1044) );
  MUX2X1 U5730 ( .B(arr[1793]), .A(arr[1826]), .S(n2466), .Y(n1038) );
  MUX2X1 U5731 ( .B(arr[1727]), .A(arr[1760]), .S(n2466), .Y(n1037) );
  MUX2X1 U5732 ( .B(arr[1661]), .A(arr[1694]), .S(n2466), .Y(n1041) );
  MUX2X1 U5733 ( .B(arr[1595]), .A(arr[1628]), .S(n2466), .Y(n1040) );
  MUX2X1 U5734 ( .B(n1039), .A(n1036), .S(n2601), .Y(n1043) );
  MUX2X1 U5735 ( .B(arr[1529]), .A(arr[1562]), .S(n2467), .Y(n1047) );
  MUX2X1 U5736 ( .B(arr[1463]), .A(arr[1496]), .S(n2467), .Y(n1046) );
  MUX2X1 U5737 ( .B(arr[1397]), .A(arr[1430]), .S(n2467), .Y(n1050) );
  MUX2X1 U5738 ( .B(arr[1331]), .A(arr[1364]), .S(n2467), .Y(n1049) );
  MUX2X1 U5739 ( .B(n1048), .A(n1045), .S(n2601), .Y(n1059) );
  MUX2X1 U5740 ( .B(arr[1265]), .A(arr[1298]), .S(n2467), .Y(n1053) );
  MUX2X1 U5741 ( .B(arr[1199]), .A(arr[1232]), .S(n2467), .Y(n1052) );
  MUX2X1 U5742 ( .B(arr[1133]), .A(arr[1166]), .S(n2467), .Y(n1056) );
  MUX2X1 U5743 ( .B(arr[1067]), .A(arr[1100]), .S(n2467), .Y(n1055) );
  MUX2X1 U5744 ( .B(n1054), .A(n1051), .S(n2601), .Y(n1058) );
  MUX2X1 U5745 ( .B(n1057), .A(n1042), .S(n2637), .Y(n1091) );
  MUX2X1 U5746 ( .B(arr[1001]), .A(arr[1034]), .S(n2467), .Y(n1062) );
  MUX2X1 U5747 ( .B(arr[935]), .A(arr[968]), .S(n2467), .Y(n1061) );
  MUX2X1 U5748 ( .B(arr[869]), .A(arr[902]), .S(n2467), .Y(n1065) );
  MUX2X1 U5749 ( .B(arr[803]), .A(arr[836]), .S(n2467), .Y(n1064) );
  MUX2X1 U5750 ( .B(n1063), .A(n1060), .S(n2601), .Y(n1074) );
  MUX2X1 U5751 ( .B(arr[737]), .A(arr[770]), .S(n2468), .Y(n1068) );
  MUX2X1 U5752 ( .B(arr[671]), .A(arr[704]), .S(n2468), .Y(n1067) );
  MUX2X1 U5753 ( .B(arr[605]), .A(arr[638]), .S(n2468), .Y(n1071) );
  MUX2X1 U5754 ( .B(arr[539]), .A(arr[572]), .S(n2468), .Y(n1070) );
  MUX2X1 U5755 ( .B(n1069), .A(n1066), .S(n2601), .Y(n1073) );
  MUX2X1 U5756 ( .B(arr[473]), .A(arr[506]), .S(n2468), .Y(n1077) );
  MUX2X1 U5757 ( .B(arr[407]), .A(arr[440]), .S(n2468), .Y(n1076) );
  MUX2X1 U5758 ( .B(arr[341]), .A(arr[374]), .S(n2468), .Y(n1080) );
  MUX2X1 U5759 ( .B(arr[275]), .A(arr[308]), .S(n2468), .Y(n1079) );
  MUX2X1 U5760 ( .B(n1078), .A(n1075), .S(n2601), .Y(n1089) );
  MUX2X1 U5761 ( .B(arr[209]), .A(arr[242]), .S(n2468), .Y(n1083) );
  MUX2X1 U5762 ( .B(arr[143]), .A(arr[176]), .S(n2468), .Y(n1082) );
  MUX2X1 U5763 ( .B(arr[77]), .A(arr[110]), .S(n2468), .Y(n1086) );
  MUX2X1 U5764 ( .B(arr[11]), .A(arr[44]), .S(n2468), .Y(n1085) );
  MUX2X1 U5765 ( .B(n1084), .A(n1081), .S(n2601), .Y(n1088) );
  MUX2X1 U5766 ( .B(n1087), .A(n1072), .S(n2637), .Y(n1090) );
  MUX2X1 U5767 ( .B(arr[2058]), .A(arr[2091]), .S(n2469), .Y(n1094) );
  MUX2X1 U5768 ( .B(arr[1992]), .A(arr[2025]), .S(n2469), .Y(n1093) );
  MUX2X1 U5769 ( .B(arr[1926]), .A(arr[1959]), .S(n2469), .Y(n1097) );
  MUX2X1 U5770 ( .B(arr[1860]), .A(arr[1893]), .S(n2469), .Y(n1096) );
  MUX2X1 U5771 ( .B(n1095), .A(n1092), .S(n2602), .Y(n1106) );
  MUX2X1 U5772 ( .B(arr[1794]), .A(arr[1827]), .S(n2469), .Y(n1100) );
  MUX2X1 U5773 ( .B(arr[1728]), .A(arr[1761]), .S(n2469), .Y(n1099) );
  MUX2X1 U5774 ( .B(arr[1662]), .A(arr[1695]), .S(n2469), .Y(n1103) );
  MUX2X1 U5775 ( .B(arr[1596]), .A(arr[1629]), .S(n2469), .Y(n1102) );
  MUX2X1 U5776 ( .B(n1101), .A(n1098), .S(n2602), .Y(n1105) );
  MUX2X1 U5777 ( .B(arr[1530]), .A(arr[1563]), .S(n2469), .Y(n1109) );
  MUX2X1 U5778 ( .B(arr[1464]), .A(arr[1497]), .S(n2469), .Y(n1108) );
  MUX2X1 U5779 ( .B(arr[1398]), .A(arr[1431]), .S(n2469), .Y(n1112) );
  MUX2X1 U5780 ( .B(arr[1332]), .A(arr[1365]), .S(n2469), .Y(n1111) );
  MUX2X1 U5781 ( .B(n1110), .A(n1107), .S(n2602), .Y(n1121) );
  MUX2X1 U5782 ( .B(arr[1266]), .A(arr[1299]), .S(n2470), .Y(n1115) );
  MUX2X1 U5783 ( .B(arr[1200]), .A(arr[1233]), .S(n2470), .Y(n1114) );
  MUX2X1 U5784 ( .B(arr[1134]), .A(arr[1167]), .S(n2470), .Y(n1118) );
  MUX2X1 U5785 ( .B(arr[1068]), .A(arr[1101]), .S(n2470), .Y(n1117) );
  MUX2X1 U5786 ( .B(n1116), .A(n1113), .S(n2602), .Y(n1120) );
  MUX2X1 U5787 ( .B(n1119), .A(n1104), .S(n2637), .Y(n1153) );
  MUX2X1 U5788 ( .B(arr[1002]), .A(arr[1035]), .S(n2470), .Y(n1124) );
  MUX2X1 U5789 ( .B(arr[936]), .A(arr[969]), .S(n2470), .Y(n1123) );
  MUX2X1 U5790 ( .B(arr[870]), .A(arr[903]), .S(n2470), .Y(n1127) );
  MUX2X1 U5791 ( .B(arr[804]), .A(arr[837]), .S(n2470), .Y(n1126) );
  MUX2X1 U5792 ( .B(n1125), .A(n1122), .S(n2602), .Y(n1136) );
  MUX2X1 U5793 ( .B(arr[738]), .A(arr[771]), .S(n2470), .Y(n1130) );
  MUX2X1 U5794 ( .B(arr[672]), .A(arr[705]), .S(n2470), .Y(n1129) );
  MUX2X1 U5795 ( .B(arr[606]), .A(arr[639]), .S(n2470), .Y(n1133) );
  MUX2X1 U5796 ( .B(arr[540]), .A(arr[573]), .S(n2470), .Y(n1132) );
  MUX2X1 U5797 ( .B(n1131), .A(n1128), .S(n2602), .Y(n1135) );
  MUX2X1 U5798 ( .B(arr[474]), .A(arr[507]), .S(n2471), .Y(n1139) );
  MUX2X1 U5799 ( .B(arr[408]), .A(arr[441]), .S(n2471), .Y(n1138) );
  MUX2X1 U5800 ( .B(arr[342]), .A(arr[375]), .S(n2471), .Y(n1142) );
  MUX2X1 U5801 ( .B(arr[276]), .A(arr[309]), .S(n2471), .Y(n1141) );
  MUX2X1 U5802 ( .B(n1140), .A(n1137), .S(n2602), .Y(n1151) );
  MUX2X1 U5803 ( .B(arr[210]), .A(arr[243]), .S(n2471), .Y(n1145) );
  MUX2X1 U5804 ( .B(arr[144]), .A(arr[177]), .S(n2471), .Y(n1144) );
  MUX2X1 U5805 ( .B(arr[78]), .A(arr[111]), .S(n2471), .Y(n1148) );
  MUX2X1 U5806 ( .B(arr[12]), .A(arr[45]), .S(n2471), .Y(n1147) );
  MUX2X1 U5807 ( .B(n1146), .A(n1143), .S(n2602), .Y(n1150) );
  MUX2X1 U5808 ( .B(n1149), .A(n1134), .S(n2637), .Y(n1152) );
  MUX2X1 U5809 ( .B(arr[2059]), .A(arr[2092]), .S(n2471), .Y(n1156) );
  MUX2X1 U5810 ( .B(arr[1993]), .A(arr[2026]), .S(n2471), .Y(n1155) );
  MUX2X1 U5811 ( .B(arr[1927]), .A(arr[1960]), .S(n2471), .Y(n1159) );
  MUX2X1 U5812 ( .B(arr[1861]), .A(arr[1894]), .S(n2471), .Y(n1158) );
  MUX2X1 U5813 ( .B(n1157), .A(n1154), .S(n2602), .Y(n1168) );
  MUX2X1 U5814 ( .B(arr[1795]), .A(arr[1828]), .S(n2472), .Y(n1162) );
  MUX2X1 U5815 ( .B(arr[1729]), .A(arr[1762]), .S(n2472), .Y(n1161) );
  MUX2X1 U5816 ( .B(arr[1663]), .A(arr[1696]), .S(n2472), .Y(n1165) );
  MUX2X1 U5817 ( .B(arr[1597]), .A(arr[1630]), .S(n2472), .Y(n1164) );
  MUX2X1 U5818 ( .B(n1163), .A(n1160), .S(n2602), .Y(n1167) );
  MUX2X1 U5819 ( .B(arr[1531]), .A(arr[1564]), .S(n2472), .Y(n1171) );
  MUX2X1 U5820 ( .B(arr[1465]), .A(arr[1498]), .S(n2472), .Y(n1170) );
  MUX2X1 U5821 ( .B(arr[1399]), .A(arr[1432]), .S(n2472), .Y(n1174) );
  MUX2X1 U5822 ( .B(arr[1333]), .A(arr[1366]), .S(n2472), .Y(n1173) );
  MUX2X1 U5823 ( .B(n1172), .A(n1169), .S(n2602), .Y(n1183) );
  MUX2X1 U5824 ( .B(arr[1267]), .A(arr[1300]), .S(n2472), .Y(n1177) );
  MUX2X1 U5825 ( .B(arr[1201]), .A(arr[1234]), .S(n2472), .Y(n1176) );
  MUX2X1 U5826 ( .B(arr[1135]), .A(arr[1168]), .S(n2472), .Y(n1180) );
  MUX2X1 U5827 ( .B(arr[1069]), .A(arr[1102]), .S(n2472), .Y(n1179) );
  MUX2X1 U5828 ( .B(n1178), .A(n1175), .S(n2602), .Y(n1182) );
  MUX2X1 U5829 ( .B(n1181), .A(n1166), .S(n2637), .Y(n1215) );
  MUX2X1 U5830 ( .B(arr[1003]), .A(arr[1036]), .S(n2473), .Y(n1186) );
  MUX2X1 U5831 ( .B(arr[937]), .A(arr[970]), .S(n2473), .Y(n1185) );
  MUX2X1 U5832 ( .B(arr[871]), .A(arr[904]), .S(n2473), .Y(n1189) );
  MUX2X1 U5833 ( .B(arr[805]), .A(arr[838]), .S(n2473), .Y(n1188) );
  MUX2X1 U5834 ( .B(n1187), .A(n1184), .S(n2603), .Y(n1198) );
  MUX2X1 U5835 ( .B(arr[739]), .A(arr[772]), .S(n2473), .Y(n1192) );
  MUX2X1 U5836 ( .B(arr[673]), .A(arr[706]), .S(n2473), .Y(n1191) );
  MUX2X1 U5837 ( .B(arr[607]), .A(arr[640]), .S(n2473), .Y(n1195) );
  MUX2X1 U5838 ( .B(arr[541]), .A(arr[574]), .S(n2473), .Y(n1194) );
  MUX2X1 U5839 ( .B(n1193), .A(n1190), .S(n2603), .Y(n1197) );
  MUX2X1 U5840 ( .B(arr[475]), .A(arr[508]), .S(n2473), .Y(n1201) );
  MUX2X1 U5841 ( .B(arr[409]), .A(arr[442]), .S(n2473), .Y(n1200) );
  MUX2X1 U5842 ( .B(arr[343]), .A(arr[376]), .S(n2473), .Y(n1204) );
  MUX2X1 U5843 ( .B(arr[277]), .A(arr[310]), .S(n2473), .Y(n1203) );
  MUX2X1 U5844 ( .B(n1202), .A(n1199), .S(n2603), .Y(n1213) );
  MUX2X1 U5845 ( .B(arr[211]), .A(arr[244]), .S(n2474), .Y(n1207) );
  MUX2X1 U5846 ( .B(arr[145]), .A(arr[178]), .S(n2474), .Y(n1206) );
  MUX2X1 U5847 ( .B(arr[79]), .A(arr[112]), .S(n2474), .Y(n1210) );
  MUX2X1 U5848 ( .B(arr[13]), .A(arr[46]), .S(n2474), .Y(n1209) );
  MUX2X1 U5849 ( .B(n1208), .A(n1205), .S(n2603), .Y(n1212) );
  MUX2X1 U5850 ( .B(n1211), .A(n1196), .S(n2637), .Y(n1214) );
  MUX2X1 U5851 ( .B(arr[2060]), .A(arr[2093]), .S(n2474), .Y(n1218) );
  MUX2X1 U5852 ( .B(arr[1994]), .A(arr[2027]), .S(n2474), .Y(n1217) );
  MUX2X1 U5853 ( .B(arr[1928]), .A(arr[1961]), .S(n2474), .Y(n1221) );
  MUX2X1 U5854 ( .B(arr[1862]), .A(arr[1895]), .S(n2474), .Y(n1220) );
  MUX2X1 U5855 ( .B(n1219), .A(n1216), .S(n2603), .Y(n1230) );
  MUX2X1 U5856 ( .B(arr[1796]), .A(arr[1829]), .S(n2474), .Y(n1224) );
  MUX2X1 U5857 ( .B(arr[1730]), .A(arr[1763]), .S(n2474), .Y(n1223) );
  MUX2X1 U5858 ( .B(arr[1664]), .A(arr[1697]), .S(n2474), .Y(n1227) );
  MUX2X1 U5859 ( .B(arr[1598]), .A(arr[1631]), .S(n2474), .Y(n1226) );
  MUX2X1 U5860 ( .B(n1225), .A(n1222), .S(n2603), .Y(n1229) );
  MUX2X1 U5861 ( .B(arr[1532]), .A(arr[1565]), .S(n2475), .Y(n1233) );
  MUX2X1 U5862 ( .B(arr[1466]), .A(arr[1499]), .S(n2475), .Y(n1232) );
  MUX2X1 U5863 ( .B(arr[1400]), .A(arr[1433]), .S(n2475), .Y(n1236) );
  MUX2X1 U5864 ( .B(arr[1334]), .A(arr[1367]), .S(n2475), .Y(n1235) );
  MUX2X1 U5865 ( .B(n1234), .A(n1231), .S(n2603), .Y(n1245) );
  MUX2X1 U5866 ( .B(arr[1268]), .A(arr[1301]), .S(n2475), .Y(n1239) );
  MUX2X1 U5867 ( .B(arr[1202]), .A(arr[1235]), .S(n2475), .Y(n1238) );
  MUX2X1 U5868 ( .B(arr[1136]), .A(arr[1169]), .S(n2475), .Y(n1242) );
  MUX2X1 U5869 ( .B(arr[1070]), .A(arr[1103]), .S(n2475), .Y(n1241) );
  MUX2X1 U5870 ( .B(n1240), .A(n1237), .S(n2603), .Y(n1244) );
  MUX2X1 U5871 ( .B(n1243), .A(n1228), .S(n2637), .Y(n1277) );
  MUX2X1 U5872 ( .B(arr[1004]), .A(arr[1037]), .S(n2475), .Y(n1248) );
  MUX2X1 U5873 ( .B(arr[938]), .A(arr[971]), .S(n2475), .Y(n1247) );
  MUX2X1 U5874 ( .B(arr[872]), .A(arr[905]), .S(n2475), .Y(n1251) );
  MUX2X1 U5875 ( .B(arr[806]), .A(arr[839]), .S(n2475), .Y(n1250) );
  MUX2X1 U5876 ( .B(n1249), .A(n1246), .S(n2603), .Y(n1260) );
  MUX2X1 U5877 ( .B(arr[740]), .A(arr[773]), .S(n2476), .Y(n1254) );
  MUX2X1 U5878 ( .B(arr[674]), .A(arr[707]), .S(n2476), .Y(n1253) );
  MUX2X1 U5879 ( .B(arr[608]), .A(arr[641]), .S(n2476), .Y(n1257) );
  MUX2X1 U5880 ( .B(arr[542]), .A(arr[575]), .S(n2476), .Y(n1256) );
  MUX2X1 U5881 ( .B(n1255), .A(n1252), .S(n2603), .Y(n1259) );
  MUX2X1 U5882 ( .B(arr[476]), .A(arr[509]), .S(n2476), .Y(n1263) );
  MUX2X1 U5883 ( .B(arr[410]), .A(arr[443]), .S(n2476), .Y(n1262) );
  MUX2X1 U5884 ( .B(arr[344]), .A(arr[377]), .S(n2476), .Y(n1266) );
  MUX2X1 U5885 ( .B(arr[278]), .A(arr[311]), .S(n2476), .Y(n1265) );
  MUX2X1 U5886 ( .B(n1264), .A(n1261), .S(n2603), .Y(n1275) );
  MUX2X1 U5887 ( .B(arr[212]), .A(arr[245]), .S(n2476), .Y(n1269) );
  MUX2X1 U5888 ( .B(arr[146]), .A(arr[179]), .S(n2476), .Y(n1268) );
  MUX2X1 U5889 ( .B(arr[80]), .A(arr[113]), .S(n2476), .Y(n1272) );
  MUX2X1 U5890 ( .B(arr[14]), .A(arr[47]), .S(n2476), .Y(n1271) );
  MUX2X1 U5891 ( .B(n1270), .A(n1267), .S(n2603), .Y(n1274) );
  MUX2X1 U5892 ( .B(n1273), .A(n1258), .S(n2637), .Y(n1276) );
  MUX2X1 U5893 ( .B(arr[2061]), .A(arr[2094]), .S(n2477), .Y(n1280) );
  MUX2X1 U5894 ( .B(arr[1995]), .A(arr[2028]), .S(n2477), .Y(n1279) );
  MUX2X1 U5895 ( .B(arr[1929]), .A(arr[1962]), .S(n2477), .Y(n1283) );
  MUX2X1 U5896 ( .B(arr[1863]), .A(arr[1896]), .S(n2477), .Y(n1282) );
  MUX2X1 U5897 ( .B(n1281), .A(n1278), .S(n2604), .Y(n1292) );
  MUX2X1 U5898 ( .B(arr[1797]), .A(arr[1830]), .S(n2477), .Y(n1286) );
  MUX2X1 U5899 ( .B(arr[1731]), .A(arr[1764]), .S(n2477), .Y(n1285) );
  MUX2X1 U5900 ( .B(arr[1665]), .A(arr[1698]), .S(n2477), .Y(n1289) );
  MUX2X1 U5901 ( .B(arr[1599]), .A(arr[1632]), .S(n2477), .Y(n1288) );
  MUX2X1 U5902 ( .B(n1287), .A(n1284), .S(n2604), .Y(n1291) );
  MUX2X1 U5903 ( .B(arr[1533]), .A(arr[1566]), .S(n2477), .Y(n1295) );
  MUX2X1 U5904 ( .B(arr[1467]), .A(arr[1500]), .S(n2477), .Y(n1294) );
  MUX2X1 U5905 ( .B(arr[1401]), .A(arr[1434]), .S(n2477), .Y(n1298) );
  MUX2X1 U5906 ( .B(arr[1335]), .A(arr[1368]), .S(n2477), .Y(n1297) );
  MUX2X1 U5907 ( .B(n1296), .A(n1293), .S(n2604), .Y(n1307) );
  MUX2X1 U5908 ( .B(arr[1269]), .A(arr[1302]), .S(n2478), .Y(n1301) );
  MUX2X1 U5909 ( .B(arr[1203]), .A(arr[1236]), .S(n2478), .Y(n1300) );
  MUX2X1 U5910 ( .B(arr[1137]), .A(arr[1170]), .S(n2478), .Y(n1304) );
  MUX2X1 U5911 ( .B(arr[1071]), .A(arr[1104]), .S(n2478), .Y(n1303) );
  MUX2X1 U5912 ( .B(n1302), .A(n1299), .S(n2604), .Y(n1306) );
  MUX2X1 U5913 ( .B(n1305), .A(n1290), .S(n2638), .Y(n1339) );
  MUX2X1 U5914 ( .B(arr[1005]), .A(arr[1038]), .S(n2478), .Y(n1310) );
  MUX2X1 U5915 ( .B(arr[939]), .A(arr[972]), .S(n2478), .Y(n1309) );
  MUX2X1 U5916 ( .B(arr[873]), .A(arr[906]), .S(n2478), .Y(n1313) );
  MUX2X1 U5917 ( .B(arr[807]), .A(arr[840]), .S(n2478), .Y(n1312) );
  MUX2X1 U5918 ( .B(n1311), .A(n1308), .S(n2604), .Y(n1322) );
  MUX2X1 U5919 ( .B(arr[741]), .A(arr[774]), .S(n2478), .Y(n1316) );
  MUX2X1 U5920 ( .B(arr[675]), .A(arr[708]), .S(n2478), .Y(n1315) );
  MUX2X1 U5921 ( .B(arr[609]), .A(arr[642]), .S(n2478), .Y(n1319) );
  MUX2X1 U5922 ( .B(arr[543]), .A(arr[576]), .S(n2478), .Y(n1318) );
  MUX2X1 U5923 ( .B(n1317), .A(n1314), .S(n2604), .Y(n1321) );
  MUX2X1 U5924 ( .B(arr[477]), .A(arr[510]), .S(n2479), .Y(n1325) );
  MUX2X1 U5925 ( .B(arr[411]), .A(arr[444]), .S(n2479), .Y(n1324) );
  MUX2X1 U5926 ( .B(arr[345]), .A(arr[378]), .S(n2479), .Y(n1328) );
  MUX2X1 U5927 ( .B(arr[279]), .A(arr[312]), .S(n2479), .Y(n1327) );
  MUX2X1 U5928 ( .B(n1326), .A(n1323), .S(n2604), .Y(n1337) );
  MUX2X1 U5929 ( .B(arr[213]), .A(arr[246]), .S(n2479), .Y(n1331) );
  MUX2X1 U5930 ( .B(arr[147]), .A(arr[180]), .S(n2479), .Y(n1330) );
  MUX2X1 U5931 ( .B(arr[81]), .A(arr[114]), .S(n2479), .Y(n1334) );
  MUX2X1 U5932 ( .B(arr[15]), .A(arr[48]), .S(n2479), .Y(n1333) );
  MUX2X1 U5933 ( .B(n1332), .A(n1329), .S(n2604), .Y(n1336) );
  MUX2X1 U5934 ( .B(n1335), .A(n1320), .S(n2638), .Y(n1338) );
  MUX2X1 U5935 ( .B(arr[2062]), .A(arr[2095]), .S(n2479), .Y(n1342) );
  MUX2X1 U5936 ( .B(arr[1996]), .A(arr[2029]), .S(n2479), .Y(n1341) );
  MUX2X1 U5937 ( .B(arr[1930]), .A(arr[1963]), .S(n2479), .Y(n1345) );
  MUX2X1 U5938 ( .B(arr[1864]), .A(arr[1897]), .S(n2479), .Y(n1344) );
  MUX2X1 U5939 ( .B(n1343), .A(n1340), .S(n2604), .Y(n1354) );
  MUX2X1 U5940 ( .B(arr[1798]), .A(arr[1831]), .S(n2480), .Y(n1348) );
  MUX2X1 U5941 ( .B(arr[1732]), .A(arr[1765]), .S(n2480), .Y(n1347) );
  MUX2X1 U5942 ( .B(arr[1666]), .A(arr[1699]), .S(n2480), .Y(n1351) );
  MUX2X1 U5943 ( .B(arr[1600]), .A(arr[1633]), .S(n2480), .Y(n1350) );
  MUX2X1 U5944 ( .B(n1349), .A(n1346), .S(n2604), .Y(n1353) );
  MUX2X1 U5945 ( .B(arr[1534]), .A(arr[1567]), .S(n2480), .Y(n1357) );
  MUX2X1 U5946 ( .B(arr[1468]), .A(arr[1501]), .S(n2480), .Y(n1356) );
  MUX2X1 U5947 ( .B(arr[1402]), .A(arr[1435]), .S(n2480), .Y(n1360) );
  MUX2X1 U5948 ( .B(arr[1336]), .A(arr[1369]), .S(n2480), .Y(n1359) );
  MUX2X1 U5949 ( .B(n1358), .A(n1355), .S(n2604), .Y(n1369) );
  MUX2X1 U5950 ( .B(arr[1270]), .A(arr[1303]), .S(n2480), .Y(n1363) );
  MUX2X1 U5951 ( .B(arr[1204]), .A(arr[1237]), .S(n2480), .Y(n1362) );
  MUX2X1 U5952 ( .B(arr[1138]), .A(arr[1171]), .S(n2480), .Y(n1366) );
  MUX2X1 U5953 ( .B(arr[1072]), .A(arr[1105]), .S(n2480), .Y(n1365) );
  MUX2X1 U5954 ( .B(n1364), .A(n1361), .S(n2604), .Y(n1368) );
  MUX2X1 U5955 ( .B(n1367), .A(n1352), .S(n2638), .Y(n1401) );
  MUX2X1 U5956 ( .B(arr[1006]), .A(arr[1039]), .S(n2481), .Y(n1372) );
  MUX2X1 U5957 ( .B(arr[940]), .A(arr[973]), .S(n2481), .Y(n1371) );
  MUX2X1 U5958 ( .B(arr[874]), .A(arr[907]), .S(n2481), .Y(n1375) );
  MUX2X1 U5959 ( .B(arr[808]), .A(arr[841]), .S(n2481), .Y(n1374) );
  MUX2X1 U5960 ( .B(n1373), .A(n1370), .S(n2605), .Y(n1384) );
  MUX2X1 U5961 ( .B(arr[742]), .A(arr[775]), .S(n2481), .Y(n1378) );
  MUX2X1 U5962 ( .B(arr[676]), .A(arr[709]), .S(n2481), .Y(n1377) );
  MUX2X1 U5963 ( .B(arr[610]), .A(arr[643]), .S(n2481), .Y(n1381) );
  MUX2X1 U5964 ( .B(arr[544]), .A(arr[577]), .S(n2481), .Y(n1380) );
  MUX2X1 U5965 ( .B(n1379), .A(n1376), .S(n2605), .Y(n1383) );
  MUX2X1 U5966 ( .B(arr[478]), .A(arr[511]), .S(n2481), .Y(n1387) );
  MUX2X1 U5967 ( .B(arr[412]), .A(arr[445]), .S(n2481), .Y(n1386) );
  MUX2X1 U5968 ( .B(arr[346]), .A(arr[379]), .S(n2481), .Y(n1390) );
  MUX2X1 U5969 ( .B(arr[280]), .A(arr[313]), .S(n2481), .Y(n1389) );
  MUX2X1 U5970 ( .B(n1388), .A(n1385), .S(n2605), .Y(n1399) );
  MUX2X1 U5971 ( .B(arr[214]), .A(arr[247]), .S(n2482), .Y(n1393) );
  MUX2X1 U5972 ( .B(arr[148]), .A(arr[181]), .S(n2482), .Y(n1392) );
  MUX2X1 U5973 ( .B(arr[82]), .A(arr[115]), .S(n2482), .Y(n1396) );
  MUX2X1 U5974 ( .B(arr[16]), .A(arr[49]), .S(n2482), .Y(n1395) );
  MUX2X1 U5975 ( .B(n1394), .A(n1391), .S(n2605), .Y(n1398) );
  MUX2X1 U5976 ( .B(n1397), .A(n1382), .S(n2638), .Y(n1400) );
  MUX2X1 U5977 ( .B(arr[2063]), .A(arr[2096]), .S(n2482), .Y(n1404) );
  MUX2X1 U5978 ( .B(arr[1997]), .A(arr[2030]), .S(n2482), .Y(n1403) );
  MUX2X1 U5979 ( .B(arr[1931]), .A(arr[1964]), .S(n2482), .Y(n1407) );
  MUX2X1 U5980 ( .B(arr[1865]), .A(arr[1898]), .S(n2482), .Y(n1406) );
  MUX2X1 U5981 ( .B(n1405), .A(n1402), .S(n2605), .Y(n1416) );
  MUX2X1 U5982 ( .B(arr[1799]), .A(arr[1832]), .S(n2482), .Y(n1410) );
  MUX2X1 U5983 ( .B(arr[1733]), .A(arr[1766]), .S(n2482), .Y(n1409) );
  MUX2X1 U5984 ( .B(arr[1667]), .A(arr[1700]), .S(n2482), .Y(n1413) );
  MUX2X1 U5985 ( .B(arr[1601]), .A(arr[1634]), .S(n2482), .Y(n1412) );
  MUX2X1 U5986 ( .B(n1411), .A(n1408), .S(n2605), .Y(n1415) );
  MUX2X1 U5987 ( .B(arr[1535]), .A(arr[1568]), .S(n2483), .Y(n1419) );
  MUX2X1 U5988 ( .B(arr[1469]), .A(arr[1502]), .S(n2483), .Y(n1418) );
  MUX2X1 U5989 ( .B(arr[1403]), .A(arr[1436]), .S(n2483), .Y(n1422) );
  MUX2X1 U5990 ( .B(arr[1337]), .A(arr[1370]), .S(n2483), .Y(n1421) );
  MUX2X1 U5991 ( .B(n1420), .A(n1417), .S(n2605), .Y(n1431) );
  MUX2X1 U5992 ( .B(arr[1271]), .A(arr[1304]), .S(n2483), .Y(n1425) );
  MUX2X1 U5993 ( .B(arr[1205]), .A(arr[1238]), .S(n2483), .Y(n1424) );
  MUX2X1 U5994 ( .B(arr[1139]), .A(arr[1172]), .S(n2483), .Y(n1428) );
  MUX2X1 U5995 ( .B(arr[1073]), .A(arr[1106]), .S(n2483), .Y(n1427) );
  MUX2X1 U5996 ( .B(n1426), .A(n1423), .S(n2605), .Y(n1430) );
  MUX2X1 U5997 ( .B(n1429), .A(n1414), .S(n2638), .Y(n1463) );
  MUX2X1 U5998 ( .B(arr[1007]), .A(arr[1040]), .S(n2483), .Y(n1434) );
  MUX2X1 U5999 ( .B(arr[941]), .A(arr[974]), .S(n2483), .Y(n1433) );
  MUX2X1 U6000 ( .B(arr[875]), .A(arr[908]), .S(n2483), .Y(n1437) );
  MUX2X1 U6001 ( .B(arr[809]), .A(arr[842]), .S(n2483), .Y(n1436) );
  MUX2X1 U6002 ( .B(n1435), .A(n1432), .S(n2605), .Y(n1446) );
  MUX2X1 U6003 ( .B(arr[743]), .A(arr[776]), .S(n2484), .Y(n1440) );
  MUX2X1 U6004 ( .B(arr[677]), .A(arr[710]), .S(n2484), .Y(n1439) );
  MUX2X1 U6005 ( .B(arr[611]), .A(arr[644]), .S(n2484), .Y(n1443) );
  MUX2X1 U6006 ( .B(arr[545]), .A(arr[578]), .S(n2484), .Y(n1442) );
  MUX2X1 U6007 ( .B(n1441), .A(n1438), .S(n2605), .Y(n1445) );
  MUX2X1 U6008 ( .B(arr[479]), .A(arr[512]), .S(n2484), .Y(n1449) );
  MUX2X1 U6009 ( .B(arr[413]), .A(arr[446]), .S(n2484), .Y(n1448) );
  MUX2X1 U6010 ( .B(arr[347]), .A(arr[380]), .S(n2484), .Y(n1452) );
  MUX2X1 U6011 ( .B(arr[281]), .A(arr[314]), .S(n2484), .Y(n1451) );
  MUX2X1 U6012 ( .B(n1450), .A(n1447), .S(n2605), .Y(n1461) );
  MUX2X1 U6013 ( .B(arr[215]), .A(arr[248]), .S(n2484), .Y(n1455) );
  MUX2X1 U6014 ( .B(arr[149]), .A(arr[182]), .S(n2484), .Y(n1454) );
  MUX2X1 U6015 ( .B(arr[83]), .A(arr[116]), .S(n2484), .Y(n1458) );
  MUX2X1 U6016 ( .B(arr[17]), .A(arr[50]), .S(n2484), .Y(n1457) );
  MUX2X1 U6017 ( .B(n1456), .A(n1453), .S(n2605), .Y(n1460) );
  MUX2X1 U6018 ( .B(n1459), .A(n1444), .S(n2638), .Y(n1462) );
  MUX2X1 U6019 ( .B(arr[2064]), .A(arr[2097]), .S(n2485), .Y(n1466) );
  MUX2X1 U6020 ( .B(arr[1998]), .A(arr[2031]), .S(n2485), .Y(n1465) );
  MUX2X1 U6021 ( .B(arr[1932]), .A(arr[1965]), .S(n2485), .Y(n1469) );
  MUX2X1 U6022 ( .B(arr[1866]), .A(arr[1899]), .S(n2485), .Y(n1468) );
  MUX2X1 U6023 ( .B(n1467), .A(n1464), .S(n2606), .Y(n1478) );
  MUX2X1 U6024 ( .B(arr[1800]), .A(arr[1833]), .S(n2485), .Y(n1472) );
  MUX2X1 U6025 ( .B(arr[1734]), .A(arr[1767]), .S(n2485), .Y(n1471) );
  MUX2X1 U6026 ( .B(arr[1668]), .A(arr[1701]), .S(n2485), .Y(n1475) );
  MUX2X1 U6027 ( .B(arr[1602]), .A(arr[1635]), .S(n2485), .Y(n1474) );
  MUX2X1 U6028 ( .B(n1473), .A(n1470), .S(n2606), .Y(n1477) );
  MUX2X1 U6029 ( .B(arr[1536]), .A(arr[1569]), .S(n2485), .Y(n1481) );
  MUX2X1 U6030 ( .B(arr[1470]), .A(arr[1503]), .S(n2485), .Y(n1480) );
  MUX2X1 U6031 ( .B(arr[1404]), .A(arr[1437]), .S(n2485), .Y(n1484) );
  MUX2X1 U6032 ( .B(arr[1338]), .A(arr[1371]), .S(n2485), .Y(n1483) );
  MUX2X1 U6033 ( .B(n1482), .A(n1479), .S(n2606), .Y(n1493) );
  MUX2X1 U6034 ( .B(arr[1272]), .A(arr[1305]), .S(n2486), .Y(n1487) );
  MUX2X1 U6035 ( .B(arr[1206]), .A(arr[1239]), .S(n2486), .Y(n1486) );
  MUX2X1 U6036 ( .B(arr[1140]), .A(arr[1173]), .S(n2486), .Y(n1490) );
  MUX2X1 U6037 ( .B(arr[1074]), .A(arr[1107]), .S(n2486), .Y(n1489) );
  MUX2X1 U6038 ( .B(n1488), .A(n1485), .S(n2606), .Y(n1492) );
  MUX2X1 U6039 ( .B(n1491), .A(n1476), .S(n2638), .Y(n1525) );
  MUX2X1 U6040 ( .B(arr[1008]), .A(arr[1041]), .S(n2486), .Y(n1496) );
  MUX2X1 U6041 ( .B(arr[942]), .A(arr[975]), .S(n2486), .Y(n1495) );
  MUX2X1 U6042 ( .B(arr[876]), .A(arr[909]), .S(n2486), .Y(n1499) );
  MUX2X1 U6043 ( .B(arr[810]), .A(arr[843]), .S(n2486), .Y(n1498) );
  MUX2X1 U6044 ( .B(n1497), .A(n1494), .S(n2606), .Y(n1508) );
  MUX2X1 U6045 ( .B(arr[744]), .A(arr[777]), .S(n2486), .Y(n1502) );
  MUX2X1 U6046 ( .B(arr[678]), .A(arr[711]), .S(n2486), .Y(n1501) );
  MUX2X1 U6047 ( .B(arr[612]), .A(arr[645]), .S(n2486), .Y(n1505) );
  MUX2X1 U6048 ( .B(arr[546]), .A(arr[579]), .S(n2486), .Y(n1504) );
  MUX2X1 U6049 ( .B(n1503), .A(n1500), .S(n2606), .Y(n1507) );
  MUX2X1 U6050 ( .B(arr[480]), .A(arr[513]), .S(n2487), .Y(n1511) );
  MUX2X1 U6051 ( .B(arr[414]), .A(arr[447]), .S(n2487), .Y(n1510) );
  MUX2X1 U6052 ( .B(arr[348]), .A(arr[381]), .S(n2487), .Y(n1514) );
  MUX2X1 U6053 ( .B(arr[282]), .A(arr[315]), .S(n2487), .Y(n1513) );
  MUX2X1 U6054 ( .B(n1512), .A(n1509), .S(n2606), .Y(n1523) );
  MUX2X1 U6055 ( .B(arr[216]), .A(arr[249]), .S(n2487), .Y(n1517) );
  MUX2X1 U6056 ( .B(arr[150]), .A(arr[183]), .S(n2487), .Y(n1516) );
  MUX2X1 U6057 ( .B(arr[84]), .A(arr[117]), .S(n2487), .Y(n1520) );
  MUX2X1 U6058 ( .B(arr[18]), .A(arr[51]), .S(n2487), .Y(n1519) );
  MUX2X1 U6059 ( .B(n1518), .A(n1515), .S(n2606), .Y(n1522) );
  MUX2X1 U6060 ( .B(n1521), .A(n1506), .S(n2638), .Y(n1524) );
  MUX2X1 U6061 ( .B(arr[2065]), .A(arr[2098]), .S(n2487), .Y(n1528) );
  MUX2X1 U6062 ( .B(arr[1999]), .A(arr[2032]), .S(n2487), .Y(n1527) );
  MUX2X1 U6063 ( .B(arr[1933]), .A(arr[1966]), .S(n2487), .Y(n1531) );
  MUX2X1 U6064 ( .B(arr[1867]), .A(arr[1900]), .S(n2487), .Y(n1530) );
  MUX2X1 U6065 ( .B(n1529), .A(n1526), .S(n2606), .Y(n1540) );
  MUX2X1 U6066 ( .B(arr[1801]), .A(arr[1834]), .S(n2488), .Y(n1534) );
  MUX2X1 U6067 ( .B(arr[1735]), .A(arr[1768]), .S(n2488), .Y(n1533) );
  MUX2X1 U6068 ( .B(arr[1669]), .A(arr[1702]), .S(n2488), .Y(n1537) );
  MUX2X1 U6069 ( .B(arr[1603]), .A(arr[1636]), .S(n2488), .Y(n1536) );
  MUX2X1 U6070 ( .B(n1535), .A(n1532), .S(n2606), .Y(n1539) );
  MUX2X1 U6071 ( .B(arr[1537]), .A(arr[1570]), .S(n2488), .Y(n1543) );
  MUX2X1 U6072 ( .B(arr[1471]), .A(arr[1504]), .S(n2488), .Y(n1542) );
  MUX2X1 U6073 ( .B(arr[1405]), .A(arr[1438]), .S(n2488), .Y(n1546) );
  MUX2X1 U6074 ( .B(arr[1339]), .A(arr[1372]), .S(n2488), .Y(n1545) );
  MUX2X1 U6075 ( .B(n1544), .A(n1541), .S(n2606), .Y(n1555) );
  MUX2X1 U6076 ( .B(arr[1273]), .A(arr[1306]), .S(n2488), .Y(n1549) );
  MUX2X1 U6077 ( .B(arr[1207]), .A(arr[1240]), .S(n2488), .Y(n1548) );
  MUX2X1 U6078 ( .B(arr[1141]), .A(arr[1174]), .S(n2488), .Y(n1552) );
  MUX2X1 U6079 ( .B(arr[1075]), .A(arr[1108]), .S(n2488), .Y(n1551) );
  MUX2X1 U6080 ( .B(n1550), .A(n1547), .S(n2606), .Y(n1554) );
  MUX2X1 U6081 ( .B(n1553), .A(n1538), .S(n2638), .Y(n1587) );
  MUX2X1 U6082 ( .B(arr[1009]), .A(arr[1042]), .S(n2489), .Y(n1558) );
  MUX2X1 U6083 ( .B(arr[943]), .A(arr[976]), .S(n2489), .Y(n1557) );
  MUX2X1 U6084 ( .B(arr[877]), .A(arr[910]), .S(n2489), .Y(n1561) );
  MUX2X1 U6085 ( .B(arr[811]), .A(arr[844]), .S(n2489), .Y(n1560) );
  MUX2X1 U6086 ( .B(n1559), .A(n1556), .S(n2607), .Y(n1570) );
  MUX2X1 U6087 ( .B(arr[745]), .A(arr[778]), .S(n2489), .Y(n1564) );
  MUX2X1 U6088 ( .B(arr[679]), .A(arr[712]), .S(n2489), .Y(n1563) );
  MUX2X1 U6089 ( .B(arr[613]), .A(arr[646]), .S(n2489), .Y(n1567) );
  MUX2X1 U6090 ( .B(arr[547]), .A(arr[580]), .S(n2489), .Y(n1566) );
  MUX2X1 U6091 ( .B(n1565), .A(n1562), .S(n2607), .Y(n1569) );
  MUX2X1 U6092 ( .B(arr[481]), .A(arr[514]), .S(n2489), .Y(n1573) );
  MUX2X1 U6093 ( .B(arr[415]), .A(arr[448]), .S(n2489), .Y(n1572) );
  MUX2X1 U6094 ( .B(arr[349]), .A(arr[382]), .S(n2489), .Y(n1576) );
  MUX2X1 U6095 ( .B(arr[283]), .A(arr[316]), .S(n2489), .Y(n1575) );
  MUX2X1 U6096 ( .B(n1574), .A(n1571), .S(n2607), .Y(n1585) );
  MUX2X1 U6097 ( .B(arr[217]), .A(arr[250]), .S(n2490), .Y(n1579) );
  MUX2X1 U6098 ( .B(arr[151]), .A(arr[184]), .S(n2490), .Y(n1578) );
  MUX2X1 U6099 ( .B(arr[85]), .A(arr[118]), .S(n2490), .Y(n1582) );
  MUX2X1 U6100 ( .B(arr[19]), .A(arr[52]), .S(n2490), .Y(n1581) );
  MUX2X1 U6101 ( .B(n1580), .A(n1577), .S(n2607), .Y(n1584) );
  MUX2X1 U6102 ( .B(n1583), .A(n1568), .S(n2638), .Y(n1586) );
  MUX2X1 U6103 ( .B(arr[2066]), .A(arr[2099]), .S(n2490), .Y(n1590) );
  MUX2X1 U6104 ( .B(arr[2000]), .A(arr[2033]), .S(n2490), .Y(n1589) );
  MUX2X1 U6105 ( .B(arr[1934]), .A(arr[1967]), .S(n2490), .Y(n1593) );
  MUX2X1 U6106 ( .B(arr[1868]), .A(arr[1901]), .S(n2490), .Y(n1592) );
  MUX2X1 U6107 ( .B(n1591), .A(n1588), .S(n2607), .Y(n1602) );
  MUX2X1 U6108 ( .B(arr[1802]), .A(arr[1835]), .S(n2490), .Y(n1596) );
  MUX2X1 U6109 ( .B(arr[1736]), .A(arr[1769]), .S(n2490), .Y(n1595) );
  MUX2X1 U6110 ( .B(arr[1670]), .A(arr[1703]), .S(n2490), .Y(n1599) );
  MUX2X1 U6111 ( .B(arr[1604]), .A(arr[1637]), .S(n2490), .Y(n1598) );
  MUX2X1 U6112 ( .B(n1597), .A(n1594), .S(n2607), .Y(n1601) );
  MUX2X1 U6113 ( .B(arr[1538]), .A(arr[1571]), .S(n2491), .Y(n1605) );
  MUX2X1 U6114 ( .B(arr[1472]), .A(arr[1505]), .S(n2491), .Y(n1604) );
  MUX2X1 U6115 ( .B(arr[1406]), .A(arr[1439]), .S(n2491), .Y(n1608) );
  MUX2X1 U6116 ( .B(arr[1340]), .A(arr[1373]), .S(n2491), .Y(n1607) );
  MUX2X1 U6117 ( .B(n1606), .A(n1603), .S(n2607), .Y(n1617) );
  MUX2X1 U6118 ( .B(arr[1274]), .A(arr[1307]), .S(n2491), .Y(n1611) );
  MUX2X1 U6119 ( .B(arr[1208]), .A(arr[1241]), .S(n2491), .Y(n1610) );
  MUX2X1 U6120 ( .B(arr[1142]), .A(arr[1175]), .S(n2491), .Y(n1614) );
  MUX2X1 U6121 ( .B(arr[1076]), .A(arr[1109]), .S(n2491), .Y(n1613) );
  MUX2X1 U6122 ( .B(n1612), .A(n1609), .S(n2607), .Y(n1616) );
  MUX2X1 U6123 ( .B(n1615), .A(n1600), .S(n2638), .Y(n1649) );
  MUX2X1 U6124 ( .B(arr[1010]), .A(arr[1043]), .S(n2491), .Y(n1620) );
  MUX2X1 U6125 ( .B(arr[944]), .A(arr[977]), .S(n2491), .Y(n1619) );
  MUX2X1 U6126 ( .B(arr[878]), .A(arr[911]), .S(n2491), .Y(n1623) );
  MUX2X1 U6127 ( .B(arr[812]), .A(arr[845]), .S(n2491), .Y(n1622) );
  MUX2X1 U6128 ( .B(n1621), .A(n1618), .S(n2607), .Y(n1632) );
  MUX2X1 U6129 ( .B(arr[746]), .A(arr[779]), .S(n2492), .Y(n1626) );
  MUX2X1 U6130 ( .B(arr[680]), .A(arr[713]), .S(n2492), .Y(n1625) );
  MUX2X1 U6131 ( .B(arr[614]), .A(arr[647]), .S(n2492), .Y(n1629) );
  MUX2X1 U6132 ( .B(arr[548]), .A(arr[581]), .S(n2492), .Y(n1628) );
  MUX2X1 U6133 ( .B(n1627), .A(n1624), .S(n2607), .Y(n1631) );
  MUX2X1 U6134 ( .B(arr[482]), .A(arr[515]), .S(n2492), .Y(n1635) );
  MUX2X1 U6135 ( .B(arr[416]), .A(arr[449]), .S(n2492), .Y(n1634) );
  MUX2X1 U6136 ( .B(arr[350]), .A(arr[383]), .S(n2492), .Y(n1638) );
  MUX2X1 U6137 ( .B(arr[284]), .A(arr[317]), .S(n2492), .Y(n1637) );
  MUX2X1 U6138 ( .B(n1636), .A(n1633), .S(n2607), .Y(n1647) );
  MUX2X1 U6139 ( .B(arr[218]), .A(arr[251]), .S(n2492), .Y(n1641) );
  MUX2X1 U6140 ( .B(arr[152]), .A(arr[185]), .S(n2492), .Y(n1640) );
  MUX2X1 U6141 ( .B(arr[86]), .A(arr[119]), .S(n2492), .Y(n1644) );
  MUX2X1 U6142 ( .B(arr[20]), .A(arr[53]), .S(n2492), .Y(n1643) );
  MUX2X1 U6143 ( .B(n1642), .A(n1639), .S(n2607), .Y(n1646) );
  MUX2X1 U6144 ( .B(n1645), .A(n1630), .S(n2638), .Y(n1648) );
  MUX2X1 U6145 ( .B(arr[2067]), .A(arr[2100]), .S(n2493), .Y(n1652) );
  MUX2X1 U6146 ( .B(arr[2001]), .A(arr[2034]), .S(n2493), .Y(n1651) );
  MUX2X1 U6147 ( .B(arr[1935]), .A(arr[1968]), .S(n2493), .Y(n1655) );
  MUX2X1 U6148 ( .B(arr[1869]), .A(arr[1902]), .S(n2493), .Y(n1654) );
  MUX2X1 U6149 ( .B(n1653), .A(n1650), .S(n2608), .Y(n1664) );
  MUX2X1 U6150 ( .B(arr[1803]), .A(arr[1836]), .S(n2493), .Y(n1658) );
  MUX2X1 U6151 ( .B(arr[1737]), .A(arr[1770]), .S(n2493), .Y(n1657) );
  MUX2X1 U6152 ( .B(arr[1671]), .A(arr[1704]), .S(n2493), .Y(n1661) );
  MUX2X1 U6153 ( .B(arr[1605]), .A(arr[1638]), .S(n2493), .Y(n1660) );
  MUX2X1 U6154 ( .B(n1659), .A(n1656), .S(n2608), .Y(n1663) );
  MUX2X1 U6155 ( .B(arr[1539]), .A(arr[1572]), .S(n2493), .Y(n1667) );
  MUX2X1 U6156 ( .B(arr[1473]), .A(arr[1506]), .S(n2493), .Y(n1666) );
  MUX2X1 U6157 ( .B(arr[1407]), .A(arr[1440]), .S(n2493), .Y(n1670) );
  MUX2X1 U6158 ( .B(arr[1341]), .A(arr[1374]), .S(n2493), .Y(n1669) );
  MUX2X1 U6159 ( .B(n1668), .A(n1665), .S(n2608), .Y(n1679) );
  MUX2X1 U6160 ( .B(arr[1275]), .A(arr[1308]), .S(n2494), .Y(n1673) );
  MUX2X1 U6161 ( .B(arr[1209]), .A(arr[1242]), .S(n2494), .Y(n1672) );
  MUX2X1 U6162 ( .B(arr[1143]), .A(arr[1176]), .S(n2494), .Y(n1676) );
  MUX2X1 U6163 ( .B(arr[1077]), .A(arr[1110]), .S(n2494), .Y(n1675) );
  MUX2X1 U6164 ( .B(n1674), .A(n1671), .S(n2608), .Y(n1678) );
  MUX2X1 U6165 ( .B(n1677), .A(n1662), .S(n2639), .Y(n1711) );
  MUX2X1 U6166 ( .B(arr[1011]), .A(arr[1044]), .S(n2494), .Y(n1682) );
  MUX2X1 U6167 ( .B(arr[945]), .A(arr[978]), .S(n2494), .Y(n1681) );
  MUX2X1 U6168 ( .B(arr[879]), .A(arr[912]), .S(n2494), .Y(n1685) );
  MUX2X1 U6169 ( .B(arr[813]), .A(arr[846]), .S(n2494), .Y(n1684) );
  MUX2X1 U6170 ( .B(n1683), .A(n1680), .S(n2608), .Y(n1694) );
  MUX2X1 U6171 ( .B(arr[747]), .A(arr[780]), .S(n2494), .Y(n1688) );
  MUX2X1 U6172 ( .B(arr[681]), .A(arr[714]), .S(n2494), .Y(n1687) );
  MUX2X1 U6173 ( .B(arr[615]), .A(arr[648]), .S(n2494), .Y(n1691) );
  MUX2X1 U6174 ( .B(arr[549]), .A(arr[582]), .S(n2494), .Y(n1690) );
  MUX2X1 U6175 ( .B(n1689), .A(n1686), .S(n2608), .Y(n1693) );
  MUX2X1 U6176 ( .B(arr[483]), .A(arr[516]), .S(n2495), .Y(n1697) );
  MUX2X1 U6177 ( .B(arr[417]), .A(arr[450]), .S(n2495), .Y(n1696) );
  MUX2X1 U6178 ( .B(arr[351]), .A(arr[384]), .S(n2495), .Y(n1700) );
  MUX2X1 U6179 ( .B(arr[285]), .A(arr[318]), .S(n2495), .Y(n1699) );
  MUX2X1 U6180 ( .B(n1698), .A(n1695), .S(n2608), .Y(n1709) );
  MUX2X1 U6181 ( .B(arr[219]), .A(arr[252]), .S(n2495), .Y(n1703) );
  MUX2X1 U6182 ( .B(arr[153]), .A(arr[186]), .S(n2495), .Y(n1702) );
  MUX2X1 U6183 ( .B(arr[87]), .A(arr[120]), .S(n2495), .Y(n1706) );
  MUX2X1 U6184 ( .B(arr[21]), .A(arr[54]), .S(n2495), .Y(n1705) );
  MUX2X1 U6185 ( .B(n1704), .A(n1701), .S(n2608), .Y(n1708) );
  MUX2X1 U6186 ( .B(n1707), .A(n1692), .S(n2639), .Y(n1710) );
  MUX2X1 U6187 ( .B(arr[2068]), .A(arr[2101]), .S(n2495), .Y(n1714) );
  MUX2X1 U6188 ( .B(arr[2002]), .A(arr[2035]), .S(n2495), .Y(n1713) );
  MUX2X1 U6189 ( .B(arr[1936]), .A(arr[1969]), .S(n2495), .Y(n1717) );
  MUX2X1 U6190 ( .B(arr[1870]), .A(arr[1903]), .S(n2495), .Y(n1716) );
  MUX2X1 U6191 ( .B(n1715), .A(n1712), .S(n2608), .Y(n1726) );
  MUX2X1 U6192 ( .B(arr[1804]), .A(arr[1837]), .S(n2496), .Y(n1720) );
  MUX2X1 U6193 ( .B(arr[1738]), .A(arr[1771]), .S(n2496), .Y(n1719) );
  MUX2X1 U6194 ( .B(arr[1672]), .A(arr[1705]), .S(n2496), .Y(n1723) );
  MUX2X1 U6195 ( .B(arr[1606]), .A(arr[1639]), .S(n2496), .Y(n1722) );
  MUX2X1 U6196 ( .B(n1721), .A(n1718), .S(n2608), .Y(n1725) );
  MUX2X1 U6197 ( .B(arr[1540]), .A(arr[1573]), .S(n2496), .Y(n1729) );
  MUX2X1 U6198 ( .B(arr[1474]), .A(arr[1507]), .S(n2496), .Y(n1728) );
  MUX2X1 U6199 ( .B(arr[1408]), .A(arr[1441]), .S(n2496), .Y(n1732) );
  MUX2X1 U6200 ( .B(arr[1342]), .A(arr[1375]), .S(n2496), .Y(n1731) );
  MUX2X1 U6201 ( .B(n1730), .A(n1727), .S(n2608), .Y(n1741) );
  MUX2X1 U6202 ( .B(arr[1276]), .A(arr[1309]), .S(n2496), .Y(n1735) );
  MUX2X1 U6203 ( .B(arr[1210]), .A(arr[1243]), .S(n2496), .Y(n1734) );
  MUX2X1 U6204 ( .B(arr[1144]), .A(arr[1177]), .S(n2496), .Y(n1738) );
  MUX2X1 U6205 ( .B(arr[1078]), .A(arr[1111]), .S(n2496), .Y(n1737) );
  MUX2X1 U6206 ( .B(n1736), .A(n1733), .S(n2608), .Y(n1740) );
  MUX2X1 U6207 ( .B(n1739), .A(n1724), .S(n2639), .Y(n1773) );
  MUX2X1 U6208 ( .B(arr[1012]), .A(arr[1045]), .S(n2497), .Y(n1744) );
  MUX2X1 U6209 ( .B(arr[946]), .A(arr[979]), .S(n2497), .Y(n1743) );
  MUX2X1 U6210 ( .B(arr[880]), .A(arr[913]), .S(n2497), .Y(n1747) );
  MUX2X1 U6211 ( .B(arr[814]), .A(arr[847]), .S(n2497), .Y(n1746) );
  MUX2X1 U6212 ( .B(n1745), .A(n1742), .S(n2609), .Y(n1756) );
  MUX2X1 U6213 ( .B(arr[748]), .A(arr[781]), .S(n2497), .Y(n1750) );
  MUX2X1 U6214 ( .B(arr[682]), .A(arr[715]), .S(n2497), .Y(n1749) );
  MUX2X1 U6215 ( .B(arr[616]), .A(arr[649]), .S(n2497), .Y(n1753) );
  MUX2X1 U6216 ( .B(arr[550]), .A(arr[583]), .S(n2497), .Y(n1752) );
  MUX2X1 U6217 ( .B(n1751), .A(n1748), .S(n2609), .Y(n1755) );
  MUX2X1 U6218 ( .B(arr[484]), .A(arr[517]), .S(n2497), .Y(n1759) );
  MUX2X1 U6219 ( .B(arr[418]), .A(arr[451]), .S(n2497), .Y(n1758) );
  MUX2X1 U6220 ( .B(arr[352]), .A(arr[385]), .S(n2497), .Y(n1762) );
  MUX2X1 U6221 ( .B(arr[286]), .A(arr[319]), .S(n2497), .Y(n1761) );
  MUX2X1 U6222 ( .B(n1760), .A(n1757), .S(n2609), .Y(n1771) );
  MUX2X1 U6223 ( .B(arr[220]), .A(arr[253]), .S(n2498), .Y(n1765) );
  MUX2X1 U6224 ( .B(arr[154]), .A(arr[187]), .S(n2498), .Y(n1764) );
  MUX2X1 U6225 ( .B(arr[88]), .A(arr[121]), .S(n2498), .Y(n1768) );
  MUX2X1 U6226 ( .B(arr[22]), .A(arr[55]), .S(n2498), .Y(n1767) );
  MUX2X1 U6227 ( .B(n1766), .A(n1763), .S(n2609), .Y(n1770) );
  MUX2X1 U6228 ( .B(n1769), .A(n1754), .S(n2639), .Y(n1772) );
  MUX2X1 U6229 ( .B(arr[2069]), .A(arr[2102]), .S(n2498), .Y(n1776) );
  MUX2X1 U6230 ( .B(arr[2003]), .A(arr[2036]), .S(n2498), .Y(n1775) );
  MUX2X1 U6231 ( .B(arr[1937]), .A(arr[1970]), .S(n2498), .Y(n1779) );
  MUX2X1 U6232 ( .B(arr[1871]), .A(arr[1904]), .S(n2498), .Y(n1778) );
  MUX2X1 U6233 ( .B(n1777), .A(n1774), .S(n2609), .Y(n1788) );
  MUX2X1 U6234 ( .B(arr[1805]), .A(arr[1838]), .S(n2498), .Y(n1782) );
  MUX2X1 U6235 ( .B(arr[1739]), .A(arr[1772]), .S(n2498), .Y(n1781) );
  MUX2X1 U6236 ( .B(arr[1673]), .A(arr[1706]), .S(n2498), .Y(n1785) );
  MUX2X1 U6237 ( .B(arr[1607]), .A(arr[1640]), .S(n2498), .Y(n1784) );
  MUX2X1 U6238 ( .B(n1783), .A(n1780), .S(n2609), .Y(n1787) );
  MUX2X1 U6239 ( .B(arr[1541]), .A(arr[1574]), .S(n2499), .Y(n1791) );
  MUX2X1 U6240 ( .B(arr[1475]), .A(arr[1508]), .S(n2499), .Y(n1790) );
  MUX2X1 U6241 ( .B(arr[1409]), .A(arr[1442]), .S(n2499), .Y(n1794) );
  MUX2X1 U6242 ( .B(arr[1343]), .A(arr[1376]), .S(n2499), .Y(n1793) );
  MUX2X1 U6243 ( .B(n1792), .A(n1789), .S(n2609), .Y(n1803) );
  MUX2X1 U6244 ( .B(arr[1277]), .A(arr[1310]), .S(n2499), .Y(n1797) );
  MUX2X1 U6245 ( .B(arr[1211]), .A(arr[1244]), .S(n2499), .Y(n1796) );
  MUX2X1 U6246 ( .B(arr[1145]), .A(arr[1178]), .S(n2499), .Y(n1800) );
  MUX2X1 U6247 ( .B(arr[1079]), .A(arr[1112]), .S(n2499), .Y(n1799) );
  MUX2X1 U6248 ( .B(n1798), .A(n1795), .S(n2609), .Y(n1802) );
  MUX2X1 U6249 ( .B(n1801), .A(n1786), .S(n2639), .Y(n1835) );
  MUX2X1 U6250 ( .B(arr[1013]), .A(arr[1046]), .S(n2499), .Y(n1806) );
  MUX2X1 U6251 ( .B(arr[947]), .A(arr[980]), .S(n2499), .Y(n1805) );
  MUX2X1 U6252 ( .B(arr[881]), .A(arr[914]), .S(n2499), .Y(n1809) );
  MUX2X1 U6253 ( .B(arr[815]), .A(arr[848]), .S(n2499), .Y(n1808) );
  MUX2X1 U6254 ( .B(n1807), .A(n1804), .S(n2609), .Y(n1818) );
  MUX2X1 U6255 ( .B(arr[749]), .A(arr[782]), .S(n2500), .Y(n1812) );
  MUX2X1 U6256 ( .B(arr[683]), .A(arr[716]), .S(n2500), .Y(n1811) );
  MUX2X1 U6257 ( .B(arr[617]), .A(arr[650]), .S(n2500), .Y(n1815) );
  MUX2X1 U6258 ( .B(arr[551]), .A(arr[584]), .S(n2500), .Y(n1814) );
  MUX2X1 U6259 ( .B(n1813), .A(n1810), .S(n2609), .Y(n1817) );
  MUX2X1 U6260 ( .B(arr[485]), .A(arr[518]), .S(n2500), .Y(n1821) );
  MUX2X1 U6261 ( .B(arr[419]), .A(arr[452]), .S(n2500), .Y(n1820) );
  MUX2X1 U6262 ( .B(arr[353]), .A(arr[386]), .S(n2500), .Y(n1824) );
  MUX2X1 U6263 ( .B(arr[287]), .A(arr[320]), .S(n2500), .Y(n1823) );
  MUX2X1 U6264 ( .B(n1822), .A(n1819), .S(n2609), .Y(n1833) );
  MUX2X1 U6265 ( .B(arr[221]), .A(arr[254]), .S(n2500), .Y(n1827) );
  MUX2X1 U6266 ( .B(arr[155]), .A(arr[188]), .S(n2500), .Y(n1826) );
  MUX2X1 U6267 ( .B(arr[89]), .A(arr[122]), .S(n2500), .Y(n1830) );
  MUX2X1 U6268 ( .B(arr[23]), .A(arr[56]), .S(n2500), .Y(n1829) );
  MUX2X1 U6269 ( .B(n1828), .A(n1825), .S(n2609), .Y(n1832) );
  MUX2X1 U6270 ( .B(n1831), .A(n1816), .S(n2639), .Y(n1834) );
  MUX2X1 U6271 ( .B(arr[2070]), .A(arr[2103]), .S(n2501), .Y(n1838) );
  MUX2X1 U6272 ( .B(arr[2004]), .A(arr[2037]), .S(n2501), .Y(n1837) );
  MUX2X1 U6273 ( .B(arr[1938]), .A(arr[1971]), .S(n2501), .Y(n1841) );
  MUX2X1 U6274 ( .B(arr[1872]), .A(arr[1905]), .S(n2501), .Y(n1840) );
  MUX2X1 U6275 ( .B(n1839), .A(n1836), .S(n2610), .Y(n1850) );
  MUX2X1 U6276 ( .B(arr[1806]), .A(arr[1839]), .S(n2501), .Y(n1844) );
  MUX2X1 U6277 ( .B(arr[1740]), .A(arr[1773]), .S(n2501), .Y(n1843) );
  MUX2X1 U6278 ( .B(arr[1674]), .A(arr[1707]), .S(n2501), .Y(n1847) );
  MUX2X1 U6279 ( .B(arr[1608]), .A(arr[1641]), .S(n2501), .Y(n1846) );
  MUX2X1 U6280 ( .B(n1845), .A(n1842), .S(n2610), .Y(n1849) );
  MUX2X1 U6281 ( .B(arr[1542]), .A(arr[1575]), .S(n2501), .Y(n1853) );
  MUX2X1 U6282 ( .B(arr[1476]), .A(arr[1509]), .S(n2501), .Y(n1852) );
  MUX2X1 U6283 ( .B(arr[1410]), .A(arr[1443]), .S(n2501), .Y(n1856) );
  MUX2X1 U6284 ( .B(arr[1344]), .A(arr[1377]), .S(n2501), .Y(n1855) );
  MUX2X1 U6285 ( .B(n1854), .A(n1851), .S(n2610), .Y(n1865) );
  MUX2X1 U6286 ( .B(arr[1278]), .A(arr[1311]), .S(n2502), .Y(n1859) );
  MUX2X1 U6287 ( .B(arr[1212]), .A(arr[1245]), .S(n2502), .Y(n1858) );
  MUX2X1 U6288 ( .B(arr[1146]), .A(arr[1179]), .S(n2502), .Y(n1862) );
  MUX2X1 U6289 ( .B(arr[1080]), .A(arr[1113]), .S(n2502), .Y(n1861) );
  MUX2X1 U6290 ( .B(n1860), .A(n1857), .S(n2610), .Y(n1864) );
  MUX2X1 U6291 ( .B(n1863), .A(n1848), .S(n2639), .Y(n1897) );
  MUX2X1 U6292 ( .B(arr[1014]), .A(arr[1047]), .S(n2502), .Y(n1868) );
  MUX2X1 U6293 ( .B(arr[948]), .A(arr[981]), .S(n2502), .Y(n1867) );
  MUX2X1 U6294 ( .B(arr[882]), .A(arr[915]), .S(n2502), .Y(n1871) );
  MUX2X1 U6295 ( .B(arr[816]), .A(arr[849]), .S(n2502), .Y(n1870) );
  MUX2X1 U6296 ( .B(n1869), .A(n1866), .S(n2610), .Y(n1880) );
  MUX2X1 U6297 ( .B(arr[750]), .A(arr[783]), .S(n2502), .Y(n1874) );
  MUX2X1 U6298 ( .B(arr[684]), .A(arr[717]), .S(n2502), .Y(n1873) );
  MUX2X1 U6299 ( .B(arr[618]), .A(arr[651]), .S(n2502), .Y(n1877) );
  MUX2X1 U6300 ( .B(arr[552]), .A(arr[585]), .S(n2502), .Y(n1876) );
  MUX2X1 U6301 ( .B(n1875), .A(n1872), .S(n2610), .Y(n1879) );
  MUX2X1 U6302 ( .B(arr[486]), .A(arr[519]), .S(n2503), .Y(n1883) );
  MUX2X1 U6303 ( .B(arr[420]), .A(arr[453]), .S(n2503), .Y(n1882) );
  MUX2X1 U6304 ( .B(arr[354]), .A(arr[387]), .S(n2503), .Y(n1886) );
  MUX2X1 U6305 ( .B(arr[288]), .A(arr[321]), .S(n2503), .Y(n1885) );
  MUX2X1 U6306 ( .B(n1884), .A(n1881), .S(n2610), .Y(n1895) );
  MUX2X1 U6307 ( .B(arr[222]), .A(arr[255]), .S(n2503), .Y(n1889) );
  MUX2X1 U6308 ( .B(arr[156]), .A(arr[189]), .S(n2503), .Y(n1888) );
  MUX2X1 U6309 ( .B(arr[90]), .A(arr[123]), .S(n2503), .Y(n1892) );
  MUX2X1 U6310 ( .B(arr[24]), .A(arr[57]), .S(n2503), .Y(n1891) );
  MUX2X1 U6311 ( .B(n1890), .A(n1887), .S(n2610), .Y(n1894) );
  MUX2X1 U6312 ( .B(n1893), .A(n1878), .S(n2639), .Y(n1896) );
  MUX2X1 U6313 ( .B(arr[2071]), .A(arr[2104]), .S(n2503), .Y(n1900) );
  MUX2X1 U6314 ( .B(arr[2005]), .A(arr[2038]), .S(n2503), .Y(n1899) );
  MUX2X1 U6315 ( .B(arr[1939]), .A(arr[1972]), .S(n2503), .Y(n1903) );
  MUX2X1 U6316 ( .B(arr[1873]), .A(arr[1906]), .S(n2503), .Y(n1902) );
  MUX2X1 U6317 ( .B(n1901), .A(n1898), .S(n2610), .Y(n1912) );
  MUX2X1 U6318 ( .B(arr[1807]), .A(arr[1840]), .S(n2504), .Y(n1906) );
  MUX2X1 U6319 ( .B(arr[1741]), .A(arr[1774]), .S(n2504), .Y(n1905) );
  MUX2X1 U6320 ( .B(arr[1675]), .A(arr[1708]), .S(n2504), .Y(n1909) );
  MUX2X1 U6321 ( .B(arr[1609]), .A(arr[1642]), .S(n2504), .Y(n1908) );
  MUX2X1 U6322 ( .B(n1907), .A(n1904), .S(n2610), .Y(n1911) );
  MUX2X1 U6323 ( .B(arr[1543]), .A(arr[1576]), .S(n2504), .Y(n1915) );
  MUX2X1 U6324 ( .B(arr[1477]), .A(arr[1510]), .S(n2504), .Y(n1914) );
  MUX2X1 U6325 ( .B(arr[1411]), .A(arr[1444]), .S(n2504), .Y(n1918) );
  MUX2X1 U6326 ( .B(arr[1345]), .A(arr[1378]), .S(n2504), .Y(n1917) );
  MUX2X1 U6327 ( .B(n1916), .A(n1913), .S(n2610), .Y(n1927) );
  MUX2X1 U6328 ( .B(arr[1279]), .A(arr[1312]), .S(n2504), .Y(n1921) );
  MUX2X1 U6329 ( .B(arr[1213]), .A(arr[1246]), .S(n2504), .Y(n1920) );
  MUX2X1 U6330 ( .B(arr[1147]), .A(arr[1180]), .S(n2504), .Y(n1924) );
  MUX2X1 U6331 ( .B(arr[1081]), .A(arr[1114]), .S(n2504), .Y(n1923) );
  MUX2X1 U6332 ( .B(n1922), .A(n1919), .S(n2610), .Y(n1926) );
  MUX2X1 U6333 ( .B(n1925), .A(n1910), .S(n2639), .Y(n1959) );
  MUX2X1 U6334 ( .B(arr[1015]), .A(arr[1048]), .S(n2505), .Y(n1930) );
  MUX2X1 U6335 ( .B(arr[949]), .A(arr[982]), .S(n2505), .Y(n1929) );
  MUX2X1 U6336 ( .B(arr[883]), .A(arr[916]), .S(n2505), .Y(n1933) );
  MUX2X1 U6337 ( .B(arr[817]), .A(arr[850]), .S(n2505), .Y(n1932) );
  MUX2X1 U6338 ( .B(n1931), .A(n1928), .S(n2611), .Y(n1942) );
  MUX2X1 U6339 ( .B(arr[751]), .A(arr[784]), .S(n2505), .Y(n1936) );
  MUX2X1 U6340 ( .B(arr[685]), .A(arr[718]), .S(n2505), .Y(n1935) );
  MUX2X1 U6341 ( .B(arr[619]), .A(arr[652]), .S(n2505), .Y(n1939) );
  MUX2X1 U6342 ( .B(arr[553]), .A(arr[586]), .S(n2505), .Y(n1938) );
  MUX2X1 U6343 ( .B(n1937), .A(n1934), .S(n2611), .Y(n1941) );
  MUX2X1 U6344 ( .B(arr[487]), .A(arr[520]), .S(n2505), .Y(n1945) );
  MUX2X1 U6345 ( .B(arr[421]), .A(arr[454]), .S(n2505), .Y(n1944) );
  MUX2X1 U6346 ( .B(arr[355]), .A(arr[388]), .S(n2505), .Y(n1948) );
  MUX2X1 U6347 ( .B(arr[289]), .A(arr[322]), .S(n2505), .Y(n1947) );
  MUX2X1 U6348 ( .B(n1946), .A(n1943), .S(n2611), .Y(n1957) );
  MUX2X1 U6349 ( .B(arr[223]), .A(arr[256]), .S(n2506), .Y(n1951) );
  MUX2X1 U6350 ( .B(arr[157]), .A(arr[190]), .S(n2506), .Y(n1950) );
  MUX2X1 U6351 ( .B(arr[91]), .A(arr[124]), .S(n2506), .Y(n1954) );
  MUX2X1 U6352 ( .B(arr[25]), .A(arr[58]), .S(n2506), .Y(n1953) );
  MUX2X1 U6353 ( .B(n1952), .A(n1949), .S(n2611), .Y(n1956) );
  MUX2X1 U6354 ( .B(n1955), .A(n1940), .S(n2639), .Y(n1958) );
  MUX2X1 U6355 ( .B(arr[2072]), .A(arr[2105]), .S(n2506), .Y(n1962) );
  MUX2X1 U6356 ( .B(arr[2006]), .A(arr[2039]), .S(n2506), .Y(n1961) );
  MUX2X1 U6357 ( .B(arr[1940]), .A(arr[1973]), .S(n2506), .Y(n1965) );
  MUX2X1 U6358 ( .B(arr[1874]), .A(arr[1907]), .S(n2506), .Y(n1964) );
  MUX2X1 U6359 ( .B(n1963), .A(n1960), .S(n2611), .Y(n1974) );
  MUX2X1 U6360 ( .B(arr[1808]), .A(arr[1841]), .S(n2506), .Y(n1968) );
  MUX2X1 U6361 ( .B(arr[1742]), .A(arr[1775]), .S(n2506), .Y(n1967) );
  MUX2X1 U6362 ( .B(arr[1676]), .A(arr[1709]), .S(n2506), .Y(n1971) );
  MUX2X1 U6363 ( .B(arr[1610]), .A(arr[1643]), .S(n2506), .Y(n1970) );
  MUX2X1 U6364 ( .B(n1969), .A(n1966), .S(n2611), .Y(n1973) );
  MUX2X1 U6365 ( .B(arr[1544]), .A(arr[1577]), .S(n2507), .Y(n1977) );
  MUX2X1 U6366 ( .B(arr[1478]), .A(arr[1511]), .S(n2507), .Y(n1976) );
  MUX2X1 U6367 ( .B(arr[1412]), .A(arr[1445]), .S(n2507), .Y(n1980) );
  MUX2X1 U6368 ( .B(arr[1346]), .A(arr[1379]), .S(n2507), .Y(n1979) );
  MUX2X1 U6369 ( .B(n1978), .A(n1975), .S(n2611), .Y(n1989) );
  MUX2X1 U6370 ( .B(arr[1280]), .A(arr[1313]), .S(n2507), .Y(n1983) );
  MUX2X1 U6371 ( .B(arr[1214]), .A(arr[1247]), .S(n2507), .Y(n1982) );
  MUX2X1 U6372 ( .B(arr[1148]), .A(arr[1181]), .S(n2507), .Y(n1986) );
  MUX2X1 U6373 ( .B(arr[1082]), .A(arr[1115]), .S(n2507), .Y(n1985) );
  MUX2X1 U6374 ( .B(n1984), .A(n1981), .S(n2611), .Y(n1988) );
  MUX2X1 U6375 ( .B(n1987), .A(n1972), .S(n2639), .Y(n2021) );
  MUX2X1 U6376 ( .B(arr[1016]), .A(arr[1049]), .S(n2507), .Y(n1992) );
  MUX2X1 U6377 ( .B(arr[950]), .A(arr[983]), .S(n2507), .Y(n1991) );
  MUX2X1 U6378 ( .B(arr[884]), .A(arr[917]), .S(n2507), .Y(n1995) );
  MUX2X1 U6379 ( .B(arr[818]), .A(arr[851]), .S(n2507), .Y(n1994) );
  MUX2X1 U6380 ( .B(n1993), .A(n1990), .S(n2611), .Y(n2004) );
  MUX2X1 U6381 ( .B(arr[752]), .A(arr[785]), .S(n2508), .Y(n1998) );
  MUX2X1 U6382 ( .B(arr[686]), .A(arr[719]), .S(n2508), .Y(n1997) );
  MUX2X1 U6383 ( .B(arr[620]), .A(arr[653]), .S(n2508), .Y(n2001) );
  MUX2X1 U6384 ( .B(arr[554]), .A(arr[587]), .S(n2508), .Y(n2000) );
  MUX2X1 U6385 ( .B(n1999), .A(n1996), .S(n2611), .Y(n2003) );
  MUX2X1 U6386 ( .B(arr[488]), .A(arr[521]), .S(n2508), .Y(n2007) );
  MUX2X1 U6387 ( .B(arr[422]), .A(arr[455]), .S(n2508), .Y(n2006) );
  MUX2X1 U6388 ( .B(arr[356]), .A(arr[389]), .S(n2508), .Y(n2010) );
  MUX2X1 U6389 ( .B(arr[290]), .A(arr[323]), .S(n2508), .Y(n2009) );
  MUX2X1 U6390 ( .B(n2008), .A(n2005), .S(n2611), .Y(n2019) );
  MUX2X1 U6391 ( .B(arr[224]), .A(arr[257]), .S(n2508), .Y(n2013) );
  MUX2X1 U6392 ( .B(arr[158]), .A(arr[191]), .S(n2508), .Y(n2012) );
  MUX2X1 U6393 ( .B(arr[92]), .A(arr[125]), .S(n2508), .Y(n2016) );
  MUX2X1 U6394 ( .B(arr[26]), .A(arr[59]), .S(n2508), .Y(n2015) );
  MUX2X1 U6395 ( .B(n2014), .A(n2011), .S(n2611), .Y(n2018) );
  MUX2X1 U6396 ( .B(n2017), .A(n2002), .S(n2639), .Y(n2020) );
  MUX2X1 U6397 ( .B(arr[2073]), .A(arr[2106]), .S(n2509), .Y(n2024) );
  MUX2X1 U6398 ( .B(arr[2007]), .A(arr[2040]), .S(n2509), .Y(n2023) );
  MUX2X1 U6399 ( .B(arr[1941]), .A(arr[1974]), .S(n2509), .Y(n2027) );
  MUX2X1 U6400 ( .B(arr[1875]), .A(arr[1908]), .S(n2509), .Y(n2026) );
  MUX2X1 U6401 ( .B(n2025), .A(n2022), .S(n2612), .Y(n2036) );
  MUX2X1 U6402 ( .B(arr[1809]), .A(arr[1842]), .S(n2509), .Y(n2030) );
  MUX2X1 U6403 ( .B(arr[1743]), .A(arr[1776]), .S(n2509), .Y(n2029) );
  MUX2X1 U6404 ( .B(arr[1677]), .A(arr[1710]), .S(n2509), .Y(n2033) );
  MUX2X1 U6405 ( .B(arr[1611]), .A(arr[1644]), .S(n2509), .Y(n2032) );
  MUX2X1 U6406 ( .B(n2031), .A(n2028), .S(n2612), .Y(n2035) );
  MUX2X1 U6407 ( .B(arr[1545]), .A(arr[1578]), .S(n2509), .Y(n2039) );
  MUX2X1 U6408 ( .B(arr[1479]), .A(arr[1512]), .S(n2509), .Y(n2038) );
  MUX2X1 U6409 ( .B(arr[1413]), .A(arr[1446]), .S(n2509), .Y(n2042) );
  MUX2X1 U6410 ( .B(arr[1347]), .A(arr[1380]), .S(n2509), .Y(n2041) );
  MUX2X1 U6411 ( .B(n2040), .A(n2037), .S(n2612), .Y(n2051) );
  MUX2X1 U6412 ( .B(arr[1281]), .A(arr[1314]), .S(n2510), .Y(n2045) );
  MUX2X1 U6413 ( .B(arr[1215]), .A(arr[1248]), .S(n2510), .Y(n2044) );
  MUX2X1 U6414 ( .B(arr[1149]), .A(arr[1182]), .S(n2510), .Y(n2048) );
  MUX2X1 U6415 ( .B(arr[1083]), .A(arr[1116]), .S(n2510), .Y(n2047) );
  MUX2X1 U6416 ( .B(n2046), .A(n2043), .S(n2612), .Y(n2050) );
  MUX2X1 U6417 ( .B(n2049), .A(n2034), .S(n2640), .Y(n2083) );
  MUX2X1 U6418 ( .B(arr[1017]), .A(arr[1050]), .S(n2510), .Y(n2054) );
  MUX2X1 U6419 ( .B(arr[951]), .A(arr[984]), .S(n2510), .Y(n2053) );
  MUX2X1 U6420 ( .B(arr[885]), .A(arr[918]), .S(n2510), .Y(n2057) );
  MUX2X1 U6421 ( .B(arr[819]), .A(arr[852]), .S(n2510), .Y(n2056) );
  MUX2X1 U6422 ( .B(n2055), .A(n2052), .S(n2612), .Y(n2066) );
  MUX2X1 U6423 ( .B(arr[753]), .A(arr[786]), .S(n2510), .Y(n2060) );
  MUX2X1 U6424 ( .B(arr[687]), .A(arr[720]), .S(n2510), .Y(n2059) );
  MUX2X1 U6425 ( .B(arr[621]), .A(arr[654]), .S(n2510), .Y(n2063) );
  MUX2X1 U6426 ( .B(arr[555]), .A(arr[588]), .S(n2510), .Y(n2062) );
  MUX2X1 U6427 ( .B(n2061), .A(n2058), .S(n2612), .Y(n2065) );
  MUX2X1 U6428 ( .B(arr[489]), .A(arr[522]), .S(n2511), .Y(n2069) );
  MUX2X1 U6429 ( .B(arr[423]), .A(arr[456]), .S(n2511), .Y(n2068) );
  MUX2X1 U6430 ( .B(arr[357]), .A(arr[390]), .S(n2511), .Y(n2072) );
  MUX2X1 U6431 ( .B(arr[291]), .A(arr[324]), .S(n2511), .Y(n2071) );
  MUX2X1 U6432 ( .B(n2070), .A(n2067), .S(n2612), .Y(n2081) );
  MUX2X1 U6433 ( .B(arr[225]), .A(arr[258]), .S(n2511), .Y(n2075) );
  MUX2X1 U6434 ( .B(arr[159]), .A(arr[192]), .S(n2511), .Y(n2074) );
  MUX2X1 U6435 ( .B(arr[93]), .A(arr[126]), .S(n2511), .Y(n2078) );
  MUX2X1 U6436 ( .B(arr[27]), .A(arr[60]), .S(n2511), .Y(n2077) );
  MUX2X1 U6437 ( .B(n2076), .A(n2073), .S(n2612), .Y(n2080) );
  MUX2X1 U6438 ( .B(n2079), .A(n2064), .S(n2640), .Y(n2082) );
  MUX2X1 U6439 ( .B(arr[2074]), .A(arr[2107]), .S(n2511), .Y(n2086) );
  MUX2X1 U6440 ( .B(arr[2008]), .A(arr[2041]), .S(n2511), .Y(n2085) );
  MUX2X1 U6441 ( .B(arr[1942]), .A(arr[1975]), .S(n2511), .Y(n2089) );
  MUX2X1 U6442 ( .B(arr[1876]), .A(arr[1909]), .S(n2511), .Y(n2088) );
  MUX2X1 U6443 ( .B(n2087), .A(n2084), .S(n2612), .Y(n2098) );
  MUX2X1 U6444 ( .B(arr[1810]), .A(arr[1843]), .S(n2512), .Y(n2092) );
  MUX2X1 U6445 ( .B(arr[1744]), .A(arr[1777]), .S(n2512), .Y(n2091) );
  MUX2X1 U6446 ( .B(arr[1678]), .A(arr[1711]), .S(n2512), .Y(n2095) );
  MUX2X1 U6447 ( .B(arr[1612]), .A(arr[1645]), .S(n2512), .Y(n2094) );
  MUX2X1 U6448 ( .B(n2093), .A(n2090), .S(n2612), .Y(n2097) );
  MUX2X1 U6449 ( .B(arr[1546]), .A(arr[1579]), .S(n2512), .Y(n2101) );
  MUX2X1 U6450 ( .B(arr[1480]), .A(arr[1513]), .S(n2512), .Y(n2100) );
  MUX2X1 U6451 ( .B(arr[1414]), .A(arr[1447]), .S(n2512), .Y(n2104) );
  MUX2X1 U6452 ( .B(arr[1348]), .A(arr[1381]), .S(n2512), .Y(n2103) );
  MUX2X1 U6453 ( .B(n2102), .A(n2099), .S(n2612), .Y(n2113) );
  MUX2X1 U6454 ( .B(arr[1282]), .A(arr[1315]), .S(n2512), .Y(n2107) );
  MUX2X1 U6455 ( .B(arr[1216]), .A(arr[1249]), .S(n2512), .Y(n2106) );
  MUX2X1 U6456 ( .B(arr[1150]), .A(arr[1183]), .S(n2512), .Y(n2110) );
  MUX2X1 U6457 ( .B(arr[1084]), .A(arr[1117]), .S(n2512), .Y(n2109) );
  MUX2X1 U6458 ( .B(n2108), .A(n2105), .S(n2612), .Y(n2112) );
  MUX2X1 U6459 ( .B(n2111), .A(n2096), .S(n2640), .Y(n2145) );
  MUX2X1 U6460 ( .B(arr[1018]), .A(arr[1051]), .S(n2513), .Y(n2116) );
  MUX2X1 U6461 ( .B(arr[952]), .A(arr[985]), .S(n2513), .Y(n2115) );
  MUX2X1 U6462 ( .B(arr[886]), .A(arr[919]), .S(n2513), .Y(n2119) );
  MUX2X1 U6463 ( .B(arr[820]), .A(arr[853]), .S(n2513), .Y(n2118) );
  MUX2X1 U6464 ( .B(n2117), .A(n2114), .S(n2613), .Y(n2128) );
  MUX2X1 U6465 ( .B(arr[754]), .A(arr[787]), .S(n2513), .Y(n2122) );
  MUX2X1 U6466 ( .B(arr[688]), .A(arr[721]), .S(n2513), .Y(n2121) );
  MUX2X1 U6467 ( .B(arr[622]), .A(arr[655]), .S(n2513), .Y(n2125) );
  MUX2X1 U6468 ( .B(arr[556]), .A(arr[589]), .S(n2513), .Y(n2124) );
  MUX2X1 U6469 ( .B(n2123), .A(n2120), .S(n2613), .Y(n2127) );
  MUX2X1 U6470 ( .B(arr[490]), .A(arr[523]), .S(n2513), .Y(n2131) );
  MUX2X1 U6471 ( .B(arr[424]), .A(arr[457]), .S(n2513), .Y(n2130) );
  MUX2X1 U6472 ( .B(arr[358]), .A(arr[391]), .S(n2513), .Y(n2134) );
  MUX2X1 U6473 ( .B(arr[292]), .A(arr[325]), .S(n2513), .Y(n2133) );
  MUX2X1 U6474 ( .B(n2132), .A(n2129), .S(n2613), .Y(n2143) );
  MUX2X1 U6475 ( .B(arr[226]), .A(arr[259]), .S(n2514), .Y(n2137) );
  MUX2X1 U6476 ( .B(arr[160]), .A(arr[193]), .S(n2514), .Y(n2136) );
  MUX2X1 U6477 ( .B(arr[94]), .A(arr[127]), .S(n2514), .Y(n2140) );
  MUX2X1 U6478 ( .B(arr[28]), .A(arr[61]), .S(n2514), .Y(n2139) );
  MUX2X1 U6479 ( .B(n2138), .A(n2135), .S(n2613), .Y(n2142) );
  MUX2X1 U6480 ( .B(n2141), .A(n2126), .S(n2640), .Y(n2144) );
  MUX2X1 U6481 ( .B(arr[2075]), .A(arr[2108]), .S(n2514), .Y(n2148) );
  MUX2X1 U6482 ( .B(arr[2009]), .A(arr[2042]), .S(n2514), .Y(n2147) );
  MUX2X1 U6483 ( .B(arr[1943]), .A(arr[1976]), .S(n2514), .Y(n2151) );
  MUX2X1 U6484 ( .B(arr[1877]), .A(arr[1910]), .S(n2514), .Y(n2150) );
  MUX2X1 U6485 ( .B(n2149), .A(n2146), .S(n2613), .Y(n2160) );
  MUX2X1 U6486 ( .B(arr[1811]), .A(arr[1844]), .S(n2514), .Y(n2154) );
  MUX2X1 U6487 ( .B(arr[1745]), .A(arr[1778]), .S(n2514), .Y(n2153) );
  MUX2X1 U6488 ( .B(arr[1679]), .A(arr[1712]), .S(n2514), .Y(n2157) );
  MUX2X1 U6489 ( .B(arr[1613]), .A(arr[1646]), .S(n2514), .Y(n2156) );
  MUX2X1 U6490 ( .B(n2155), .A(n2152), .S(n2613), .Y(n2159) );
  MUX2X1 U6491 ( .B(arr[1547]), .A(arr[1580]), .S(n2515), .Y(n2163) );
  MUX2X1 U6492 ( .B(arr[1481]), .A(arr[1514]), .S(n2515), .Y(n2162) );
  MUX2X1 U6493 ( .B(arr[1415]), .A(arr[1448]), .S(n2515), .Y(n2166) );
  MUX2X1 U6494 ( .B(arr[1349]), .A(arr[1382]), .S(n2515), .Y(n2165) );
  MUX2X1 U6495 ( .B(n2164), .A(n2161), .S(n2613), .Y(n2175) );
  MUX2X1 U6496 ( .B(arr[1283]), .A(arr[1316]), .S(n2515), .Y(n2169) );
  MUX2X1 U6497 ( .B(arr[1217]), .A(arr[1250]), .S(n2515), .Y(n2168) );
  MUX2X1 U6498 ( .B(arr[1151]), .A(arr[1184]), .S(n2515), .Y(n2172) );
  MUX2X1 U6499 ( .B(arr[1085]), .A(arr[1118]), .S(n2515), .Y(n2171) );
  MUX2X1 U6500 ( .B(n2170), .A(n2167), .S(n2613), .Y(n2174) );
  MUX2X1 U6501 ( .B(n2173), .A(n2158), .S(n2640), .Y(n2207) );
  MUX2X1 U6502 ( .B(arr[1019]), .A(arr[1052]), .S(n2515), .Y(n2178) );
  MUX2X1 U6503 ( .B(arr[953]), .A(arr[986]), .S(n2515), .Y(n2177) );
  MUX2X1 U6504 ( .B(arr[887]), .A(arr[920]), .S(n2515), .Y(n2181) );
  MUX2X1 U6505 ( .B(arr[821]), .A(arr[854]), .S(n2515), .Y(n2180) );
  MUX2X1 U6506 ( .B(n2179), .A(n2176), .S(n2613), .Y(n2190) );
  MUX2X1 U6507 ( .B(arr[755]), .A(arr[788]), .S(n2516), .Y(n2184) );
  MUX2X1 U6508 ( .B(arr[689]), .A(arr[722]), .S(n2516), .Y(n2183) );
  MUX2X1 U6509 ( .B(arr[623]), .A(arr[656]), .S(n2516), .Y(n2187) );
  MUX2X1 U6510 ( .B(arr[557]), .A(arr[590]), .S(n2516), .Y(n2186) );
  MUX2X1 U6511 ( .B(n2185), .A(n2182), .S(n2613), .Y(n2189) );
  MUX2X1 U6512 ( .B(arr[491]), .A(arr[524]), .S(n2516), .Y(n2193) );
  MUX2X1 U6513 ( .B(arr[425]), .A(arr[458]), .S(n2516), .Y(n2192) );
  MUX2X1 U6514 ( .B(arr[359]), .A(arr[392]), .S(n2516), .Y(n2196) );
  MUX2X1 U6515 ( .B(arr[293]), .A(arr[326]), .S(n2516), .Y(n2195) );
  MUX2X1 U6516 ( .B(n2194), .A(n2191), .S(n2613), .Y(n2205) );
  MUX2X1 U6517 ( .B(arr[227]), .A(arr[260]), .S(n2516), .Y(n2199) );
  MUX2X1 U6518 ( .B(arr[161]), .A(arr[194]), .S(n2516), .Y(n2198) );
  MUX2X1 U6519 ( .B(arr[95]), .A(arr[128]), .S(n2516), .Y(n2202) );
  MUX2X1 U6520 ( .B(arr[29]), .A(arr[62]), .S(n2516), .Y(n2201) );
  MUX2X1 U6521 ( .B(n2200), .A(n2197), .S(n2613), .Y(n2204) );
  MUX2X1 U6522 ( .B(n2203), .A(n2188), .S(n2640), .Y(n2206) );
  MUX2X1 U6523 ( .B(arr[2076]), .A(arr[2109]), .S(n2517), .Y(n2210) );
  MUX2X1 U6524 ( .B(arr[2010]), .A(arr[2043]), .S(n2517), .Y(n2209) );
  MUX2X1 U6525 ( .B(arr[1944]), .A(arr[1977]), .S(n2517), .Y(n2226) );
  MUX2X1 U6526 ( .B(arr[1878]), .A(arr[1911]), .S(n2517), .Y(n2212) );
  MUX2X1 U6527 ( .B(n2211), .A(n2208), .S(n2614), .Y(n2235) );
  MUX2X1 U6528 ( .B(arr[1812]), .A(arr[1845]), .S(n2517), .Y(n2229) );
  MUX2X1 U6529 ( .B(arr[1746]), .A(arr[1779]), .S(n2517), .Y(n2228) );
  MUX2X1 U6530 ( .B(arr[1680]), .A(arr[1713]), .S(n2517), .Y(n2232) );
  MUX2X1 U6531 ( .B(arr[1614]), .A(arr[1647]), .S(n2517), .Y(n2231) );
  MUX2X1 U6532 ( .B(n2230), .A(n2227), .S(n2614), .Y(n2234) );
  MUX2X1 U6533 ( .B(arr[1548]), .A(arr[1581]), .S(n2517), .Y(n2238) );
  MUX2X1 U6534 ( .B(arr[1482]), .A(arr[1515]), .S(n2517), .Y(n2237) );
  MUX2X1 U6535 ( .B(arr[1416]), .A(arr[1449]), .S(n2517), .Y(n2241) );
  MUX2X1 U6536 ( .B(arr[1350]), .A(arr[1383]), .S(n2517), .Y(n2240) );
  MUX2X1 U6537 ( .B(n2239), .A(n2236), .S(n2614), .Y(n2250) );
  MUX2X1 U6538 ( .B(arr[1284]), .A(arr[1317]), .S(n2518), .Y(n2244) );
  MUX2X1 U6539 ( .B(arr[1218]), .A(arr[1251]), .S(n2518), .Y(n2243) );
  MUX2X1 U6540 ( .B(arr[1152]), .A(arr[1185]), .S(n2518), .Y(n2247) );
  MUX2X1 U6541 ( .B(arr[1086]), .A(arr[1119]), .S(n2518), .Y(n2246) );
  MUX2X1 U6542 ( .B(n2245), .A(n2242), .S(n2614), .Y(n2249) );
  MUX2X1 U6543 ( .B(n2248), .A(n2233), .S(n2640), .Y(n2282) );
  MUX2X1 U6544 ( .B(arr[1020]), .A(arr[1053]), .S(n2518), .Y(n2253) );
  MUX2X1 U6545 ( .B(arr[954]), .A(arr[987]), .S(n2518), .Y(n2252) );
  MUX2X1 U6546 ( .B(arr[888]), .A(arr[921]), .S(n2518), .Y(n2256) );
  MUX2X1 U6547 ( .B(arr[822]), .A(arr[855]), .S(n2518), .Y(n2255) );
  MUX2X1 U6548 ( .B(n2254), .A(n2251), .S(n2614), .Y(n2265) );
  MUX2X1 U6549 ( .B(arr[756]), .A(arr[789]), .S(n2518), .Y(n2259) );
  MUX2X1 U6550 ( .B(arr[690]), .A(arr[723]), .S(n2518), .Y(n2258) );
  MUX2X1 U6551 ( .B(arr[624]), .A(arr[657]), .S(n2518), .Y(n2262) );
  MUX2X1 U6552 ( .B(arr[558]), .A(arr[591]), .S(n2518), .Y(n2261) );
  MUX2X1 U6553 ( .B(n2260), .A(n2257), .S(n2614), .Y(n2264) );
  MUX2X1 U6554 ( .B(arr[492]), .A(arr[525]), .S(n2519), .Y(n2268) );
  MUX2X1 U6555 ( .B(arr[426]), .A(arr[459]), .S(n2519), .Y(n2267) );
  MUX2X1 U6556 ( .B(arr[360]), .A(arr[393]), .S(n2519), .Y(n2271) );
  MUX2X1 U6557 ( .B(arr[294]), .A(arr[327]), .S(n2519), .Y(n2270) );
  MUX2X1 U6558 ( .B(n2269), .A(n2266), .S(n2614), .Y(n2280) );
  MUX2X1 U6559 ( .B(arr[228]), .A(arr[261]), .S(n2519), .Y(n2274) );
  MUX2X1 U6560 ( .B(arr[162]), .A(arr[195]), .S(n2519), .Y(n2273) );
  MUX2X1 U6561 ( .B(arr[96]), .A(arr[129]), .S(n2519), .Y(n2277) );
  MUX2X1 U6562 ( .B(arr[30]), .A(arr[63]), .S(n2519), .Y(n2276) );
  MUX2X1 U6563 ( .B(n2275), .A(n2272), .S(n2614), .Y(n2279) );
  MUX2X1 U6564 ( .B(n2278), .A(n2263), .S(n2640), .Y(n2281) );
  MUX2X1 U6565 ( .B(arr[2077]), .A(arr[2110]), .S(n2519), .Y(n2285) );
  MUX2X1 U6566 ( .B(arr[2011]), .A(arr[2044]), .S(n2519), .Y(n2284) );
  MUX2X1 U6567 ( .B(arr[1945]), .A(arr[1978]), .S(n2519), .Y(n2288) );
  MUX2X1 U6568 ( .B(arr[1879]), .A(arr[1912]), .S(n2519), .Y(n2287) );
  MUX2X1 U6569 ( .B(n2286), .A(n2283), .S(n2614), .Y(n2297) );
  MUX2X1 U6570 ( .B(arr[1813]), .A(arr[1846]), .S(n2520), .Y(n2291) );
  MUX2X1 U6571 ( .B(arr[1747]), .A(arr[1780]), .S(n2520), .Y(n2290) );
  MUX2X1 U6572 ( .B(arr[1681]), .A(arr[1714]), .S(n2520), .Y(n2294) );
  MUX2X1 U6573 ( .B(arr[1615]), .A(arr[1648]), .S(n2520), .Y(n2293) );
  MUX2X1 U6574 ( .B(n2292), .A(n2289), .S(n2614), .Y(n2296) );
  MUX2X1 U6575 ( .B(arr[1549]), .A(arr[1582]), .S(n2520), .Y(n2300) );
  MUX2X1 U6576 ( .B(arr[1483]), .A(arr[1516]), .S(n2520), .Y(n2299) );
  MUX2X1 U6577 ( .B(arr[1417]), .A(arr[1450]), .S(n2520), .Y(n2303) );
  MUX2X1 U6578 ( .B(arr[1351]), .A(arr[1384]), .S(n2520), .Y(n2302) );
  MUX2X1 U6579 ( .B(n2301), .A(n2298), .S(n2614), .Y(n2312) );
  MUX2X1 U6580 ( .B(arr[1285]), .A(arr[1318]), .S(n2520), .Y(n2306) );
  MUX2X1 U6581 ( .B(arr[1219]), .A(arr[1252]), .S(n2520), .Y(n2305) );
  MUX2X1 U6582 ( .B(arr[1153]), .A(arr[1186]), .S(n2520), .Y(n2309) );
  MUX2X1 U6583 ( .B(arr[1087]), .A(arr[1120]), .S(n2520), .Y(n2308) );
  MUX2X1 U6584 ( .B(n2307), .A(n2304), .S(n2614), .Y(n2311) );
  MUX2X1 U6585 ( .B(n2310), .A(n2295), .S(n2640), .Y(n2344) );
  MUX2X1 U6586 ( .B(arr[1021]), .A(arr[1054]), .S(n2521), .Y(n2315) );
  MUX2X1 U6587 ( .B(arr[955]), .A(arr[988]), .S(n2521), .Y(n2314) );
  MUX2X1 U6588 ( .B(arr[889]), .A(arr[922]), .S(n2521), .Y(n2318) );
  MUX2X1 U6589 ( .B(arr[823]), .A(arr[856]), .S(n2521), .Y(n2317) );
  MUX2X1 U6590 ( .B(n2316), .A(n2313), .S(n2615), .Y(n2327) );
  MUX2X1 U6591 ( .B(arr[757]), .A(arr[790]), .S(n2521), .Y(n2321) );
  MUX2X1 U6592 ( .B(arr[691]), .A(arr[724]), .S(n2521), .Y(n2320) );
  MUX2X1 U6593 ( .B(arr[625]), .A(arr[658]), .S(n2521), .Y(n2324) );
  MUX2X1 U6594 ( .B(arr[559]), .A(arr[592]), .S(n2521), .Y(n2323) );
  MUX2X1 U6595 ( .B(n2322), .A(n2319), .S(n2615), .Y(n2326) );
  MUX2X1 U6596 ( .B(arr[493]), .A(arr[526]), .S(n2521), .Y(n2330) );
  MUX2X1 U6597 ( .B(arr[427]), .A(arr[460]), .S(n2521), .Y(n2329) );
  MUX2X1 U6598 ( .B(arr[361]), .A(arr[394]), .S(n2521), .Y(n2333) );
  MUX2X1 U6599 ( .B(arr[295]), .A(arr[328]), .S(n2521), .Y(n2332) );
  MUX2X1 U6600 ( .B(n2331), .A(n2328), .S(n2615), .Y(n2342) );
  MUX2X1 U6601 ( .B(arr[229]), .A(arr[262]), .S(n2522), .Y(n2336) );
  MUX2X1 U6602 ( .B(arr[163]), .A(arr[196]), .S(n2522), .Y(n2335) );
  MUX2X1 U6603 ( .B(arr[97]), .A(arr[130]), .S(n2522), .Y(n2339) );
  MUX2X1 U6604 ( .B(arr[31]), .A(arr[64]), .S(n2522), .Y(n2338) );
  MUX2X1 U6605 ( .B(n2337), .A(n2334), .S(n2615), .Y(n2341) );
  MUX2X1 U6606 ( .B(n2340), .A(n2325), .S(n2640), .Y(n2343) );
  MUX2X1 U6607 ( .B(arr[2078]), .A(arr[2111]), .S(n2522), .Y(n2347) );
  MUX2X1 U6608 ( .B(arr[2012]), .A(arr[2045]), .S(n2522), .Y(n2346) );
  MUX2X1 U6609 ( .B(arr[1946]), .A(arr[1979]), .S(n2522), .Y(n2350) );
  MUX2X1 U6610 ( .B(arr[1880]), .A(arr[1913]), .S(n2522), .Y(n2349) );
  MUX2X1 U6611 ( .B(n2348), .A(n2345), .S(n2615), .Y(n2359) );
  MUX2X1 U6612 ( .B(arr[1814]), .A(arr[1847]), .S(n2522), .Y(n2353) );
  MUX2X1 U6613 ( .B(arr[1748]), .A(arr[1781]), .S(n2522), .Y(n2352) );
  MUX2X1 U6614 ( .B(arr[1682]), .A(arr[1715]), .S(n2522), .Y(n2356) );
  MUX2X1 U6615 ( .B(arr[1616]), .A(arr[1649]), .S(n2522), .Y(n2355) );
  MUX2X1 U6616 ( .B(n2354), .A(n2351), .S(n2615), .Y(n2358) );
  MUX2X1 U6617 ( .B(arr[1550]), .A(arr[1583]), .S(n2523), .Y(n2362) );
  MUX2X1 U6618 ( .B(arr[1484]), .A(arr[1517]), .S(n2523), .Y(n2361) );
  MUX2X1 U6619 ( .B(arr[1418]), .A(arr[1451]), .S(n2523), .Y(n2365) );
  MUX2X1 U6620 ( .B(arr[1352]), .A(arr[1385]), .S(n2523), .Y(n2364) );
  MUX2X1 U6621 ( .B(n2363), .A(n2360), .S(n2615), .Y(n2374) );
  MUX2X1 U6622 ( .B(arr[1286]), .A(arr[1319]), .S(n2523), .Y(n2368) );
  MUX2X1 U6623 ( .B(arr[1220]), .A(arr[1253]), .S(n2523), .Y(n2367) );
  MUX2X1 U6624 ( .B(arr[1154]), .A(arr[1187]), .S(n2523), .Y(n2371) );
  MUX2X1 U6625 ( .B(arr[1088]), .A(arr[1121]), .S(n2523), .Y(n2370) );
  MUX2X1 U6626 ( .B(n2369), .A(n2366), .S(n2615), .Y(n2373) );
  MUX2X1 U6627 ( .B(n2372), .A(n2357), .S(n2640), .Y(n2406) );
  MUX2X1 U6628 ( .B(arr[1022]), .A(arr[1055]), .S(n2523), .Y(n2377) );
  MUX2X1 U6629 ( .B(arr[956]), .A(arr[989]), .S(n2523), .Y(n2376) );
  MUX2X1 U6630 ( .B(arr[890]), .A(arr[923]), .S(n2523), .Y(n2380) );
  MUX2X1 U6631 ( .B(arr[824]), .A(arr[857]), .S(n2523), .Y(n2379) );
  MUX2X1 U6632 ( .B(n2378), .A(n2375), .S(n2615), .Y(n2389) );
  MUX2X1 U6633 ( .B(arr[758]), .A(arr[791]), .S(n2524), .Y(n2383) );
  MUX2X1 U6634 ( .B(arr[692]), .A(arr[725]), .S(n2524), .Y(n2382) );
  MUX2X1 U6635 ( .B(arr[626]), .A(arr[659]), .S(n2524), .Y(n2386) );
  MUX2X1 U6636 ( .B(arr[560]), .A(arr[593]), .S(n2524), .Y(n2385) );
  MUX2X1 U6637 ( .B(n2384), .A(n2381), .S(n2615), .Y(n2388) );
  MUX2X1 U6638 ( .B(arr[494]), .A(arr[527]), .S(n2524), .Y(n2392) );
  MUX2X1 U6639 ( .B(arr[428]), .A(arr[461]), .S(n2524), .Y(n2391) );
  MUX2X1 U6640 ( .B(arr[362]), .A(arr[395]), .S(n2524), .Y(n2395) );
  MUX2X1 U6641 ( .B(arr[296]), .A(arr[329]), .S(n2524), .Y(n2394) );
  MUX2X1 U6642 ( .B(n2393), .A(n2390), .S(n2615), .Y(n2404) );
  MUX2X1 U6643 ( .B(arr[230]), .A(arr[263]), .S(n2524), .Y(n2398) );
  MUX2X1 U6644 ( .B(arr[164]), .A(arr[197]), .S(n2524), .Y(n2397) );
  MUX2X1 U6645 ( .B(arr[98]), .A(arr[131]), .S(n2524), .Y(n2401) );
  MUX2X1 U6646 ( .B(arr[32]), .A(arr[65]), .S(n2524), .Y(n2400) );
  MUX2X1 U6647 ( .B(n2399), .A(n2396), .S(n2615), .Y(n2403) );
  MUX2X1 U6648 ( .B(n2402), .A(n2387), .S(n2640), .Y(n2405) );
  AND2X2 U6649 ( .A(n6721), .B(n6720), .Y(n5607) );
  INVX1 U6650 ( .A(n6721), .Y(n6719) );
  INVX1 U6651 ( .A(fillcount[5]), .Y(n6723) );
  AND2X2 U6652 ( .A(n6677), .B(wr_ptr[0]), .Y(n5678) );
  AND2X2 U6653 ( .A(n6677), .B(n5572), .Y(n5643) );
  AND2X2 U6654 ( .A(wr_ptr[0]), .B(n5571), .Y(n4569) );
  AND2X2 U6655 ( .A(n5571), .B(n5572), .Y(n4533) );
endmodule


module FIFO_DEPTH_P26_WIDTH16 ( clk, reset, data_in, put, get, data_out, empty, 
        full, fillcount );
  input [15:0] data_in;
  output [15:0] data_out;
  output [6:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   n13, n14, n15, n16, n17, n18, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337;
  wire   [5:0] wr_ptr;
  wire   [1023:0] arr;

  DFFPOSX1 fillcount_reg_0_ ( .D(n4513), .CLK(clk), .Q(fillcount[0]) );
  DFFPOSX1 fillcount_reg_1_ ( .D(n4512), .CLK(clk), .Q(fillcount[1]) );
  DFFPOSX1 fillcount_reg_6_ ( .D(n4511), .CLK(clk), .Q(fillcount[6]) );
  DFFPOSX1 fillcount_reg_2_ ( .D(n4510), .CLK(clk), .Q(fillcount[2]) );
  DFFPOSX1 fillcount_reg_3_ ( .D(n4509), .CLK(clk), .Q(fillcount[3]) );
  DFFPOSX1 fillcount_reg_4_ ( .D(n4508), .CLK(clk), .Q(fillcount[4]) );
  DFFPOSX1 fillcount_reg_5_ ( .D(n4507), .CLK(clk), .Q(fillcount[5]) );
  DFFPOSX1 wr_ptr_reg_0_ ( .D(n4506), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n4505), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n4504), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n4503), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n4502), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 wr_ptr_reg_5_ ( .D(n4501), .CLK(clk), .Q(wr_ptr[5]) );
  DFFPOSX1 arr_reg_63__15_ ( .D(n4500), .CLK(clk), .Q(arr[1023]) );
  DFFPOSX1 arr_reg_63__14_ ( .D(n4499), .CLK(clk), .Q(arr[1022]) );
  DFFPOSX1 arr_reg_63__13_ ( .D(n4498), .CLK(clk), .Q(arr[1021]) );
  DFFPOSX1 arr_reg_63__12_ ( .D(n4497), .CLK(clk), .Q(arr[1020]) );
  DFFPOSX1 arr_reg_63__11_ ( .D(n4496), .CLK(clk), .Q(arr[1019]) );
  DFFPOSX1 arr_reg_63__10_ ( .D(n4495), .CLK(clk), .Q(arr[1018]) );
  DFFPOSX1 arr_reg_63__9_ ( .D(n4494), .CLK(clk), .Q(arr[1017]) );
  DFFPOSX1 arr_reg_63__8_ ( .D(n4493), .CLK(clk), .Q(arr[1016]) );
  DFFPOSX1 arr_reg_63__7_ ( .D(n4492), .CLK(clk), .Q(arr[1015]) );
  DFFPOSX1 arr_reg_63__6_ ( .D(n4491), .CLK(clk), .Q(arr[1014]) );
  DFFPOSX1 arr_reg_63__5_ ( .D(n4490), .CLK(clk), .Q(arr[1013]) );
  DFFPOSX1 arr_reg_63__4_ ( .D(n4489), .CLK(clk), .Q(arr[1012]) );
  DFFPOSX1 arr_reg_63__3_ ( .D(n4488), .CLK(clk), .Q(arr[1011]) );
  DFFPOSX1 arr_reg_63__2_ ( .D(n4487), .CLK(clk), .Q(arr[1010]) );
  DFFPOSX1 arr_reg_63__1_ ( .D(n4486), .CLK(clk), .Q(arr[1009]) );
  DFFPOSX1 arr_reg_63__0_ ( .D(n4485), .CLK(clk), .Q(arr[1008]) );
  DFFPOSX1 arr_reg_62__15_ ( .D(n4484), .CLK(clk), .Q(arr[1007]) );
  DFFPOSX1 arr_reg_62__14_ ( .D(n4483), .CLK(clk), .Q(arr[1006]) );
  DFFPOSX1 arr_reg_62__13_ ( .D(n4482), .CLK(clk), .Q(arr[1005]) );
  DFFPOSX1 arr_reg_62__12_ ( .D(n4481), .CLK(clk), .Q(arr[1004]) );
  DFFPOSX1 arr_reg_62__11_ ( .D(n4480), .CLK(clk), .Q(arr[1003]) );
  DFFPOSX1 arr_reg_62__10_ ( .D(n4479), .CLK(clk), .Q(arr[1002]) );
  DFFPOSX1 arr_reg_62__9_ ( .D(n4478), .CLK(clk), .Q(arr[1001]) );
  DFFPOSX1 arr_reg_62__8_ ( .D(n4477), .CLK(clk), .Q(arr[1000]) );
  DFFPOSX1 arr_reg_62__7_ ( .D(n4476), .CLK(clk), .Q(arr[999]) );
  DFFPOSX1 arr_reg_62__6_ ( .D(n4475), .CLK(clk), .Q(arr[998]) );
  DFFPOSX1 arr_reg_62__5_ ( .D(n4474), .CLK(clk), .Q(arr[997]) );
  DFFPOSX1 arr_reg_62__4_ ( .D(n4473), .CLK(clk), .Q(arr[996]) );
  DFFPOSX1 arr_reg_62__3_ ( .D(n4472), .CLK(clk), .Q(arr[995]) );
  DFFPOSX1 arr_reg_62__2_ ( .D(n4471), .CLK(clk), .Q(arr[994]) );
  DFFPOSX1 arr_reg_62__1_ ( .D(n4470), .CLK(clk), .Q(arr[993]) );
  DFFPOSX1 arr_reg_62__0_ ( .D(n4469), .CLK(clk), .Q(arr[992]) );
  DFFPOSX1 arr_reg_61__15_ ( .D(n4468), .CLK(clk), .Q(arr[991]) );
  DFFPOSX1 arr_reg_61__14_ ( .D(n4467), .CLK(clk), .Q(arr[990]) );
  DFFPOSX1 arr_reg_61__13_ ( .D(n4466), .CLK(clk), .Q(arr[989]) );
  DFFPOSX1 arr_reg_61__12_ ( .D(n4465), .CLK(clk), .Q(arr[988]) );
  DFFPOSX1 arr_reg_61__11_ ( .D(n4464), .CLK(clk), .Q(arr[987]) );
  DFFPOSX1 arr_reg_61__10_ ( .D(n4463), .CLK(clk), .Q(arr[986]) );
  DFFPOSX1 arr_reg_61__9_ ( .D(n4462), .CLK(clk), .Q(arr[985]) );
  DFFPOSX1 arr_reg_61__8_ ( .D(n4461), .CLK(clk), .Q(arr[984]) );
  DFFPOSX1 arr_reg_61__7_ ( .D(n4460), .CLK(clk), .Q(arr[983]) );
  DFFPOSX1 arr_reg_61__6_ ( .D(n4459), .CLK(clk), .Q(arr[982]) );
  DFFPOSX1 arr_reg_61__5_ ( .D(n4458), .CLK(clk), .Q(arr[981]) );
  DFFPOSX1 arr_reg_61__4_ ( .D(n4457), .CLK(clk), .Q(arr[980]) );
  DFFPOSX1 arr_reg_61__3_ ( .D(n4456), .CLK(clk), .Q(arr[979]) );
  DFFPOSX1 arr_reg_61__2_ ( .D(n4455), .CLK(clk), .Q(arr[978]) );
  DFFPOSX1 arr_reg_61__1_ ( .D(n4454), .CLK(clk), .Q(arr[977]) );
  DFFPOSX1 arr_reg_61__0_ ( .D(n4453), .CLK(clk), .Q(arr[976]) );
  DFFPOSX1 arr_reg_60__15_ ( .D(n4452), .CLK(clk), .Q(arr[975]) );
  DFFPOSX1 arr_reg_60__14_ ( .D(n4451), .CLK(clk), .Q(arr[974]) );
  DFFPOSX1 arr_reg_60__13_ ( .D(n4450), .CLK(clk), .Q(arr[973]) );
  DFFPOSX1 arr_reg_60__12_ ( .D(n4449), .CLK(clk), .Q(arr[972]) );
  DFFPOSX1 arr_reg_60__11_ ( .D(n4448), .CLK(clk), .Q(arr[971]) );
  DFFPOSX1 arr_reg_60__10_ ( .D(n4447), .CLK(clk), .Q(arr[970]) );
  DFFPOSX1 arr_reg_60__9_ ( .D(n4446), .CLK(clk), .Q(arr[969]) );
  DFFPOSX1 arr_reg_60__8_ ( .D(n4445), .CLK(clk), .Q(arr[968]) );
  DFFPOSX1 arr_reg_60__7_ ( .D(n4444), .CLK(clk), .Q(arr[967]) );
  DFFPOSX1 arr_reg_60__6_ ( .D(n4443), .CLK(clk), .Q(arr[966]) );
  DFFPOSX1 arr_reg_60__5_ ( .D(n4442), .CLK(clk), .Q(arr[965]) );
  DFFPOSX1 arr_reg_60__4_ ( .D(n4441), .CLK(clk), .Q(arr[964]) );
  DFFPOSX1 arr_reg_60__3_ ( .D(n4440), .CLK(clk), .Q(arr[963]) );
  DFFPOSX1 arr_reg_60__2_ ( .D(n4439), .CLK(clk), .Q(arr[962]) );
  DFFPOSX1 arr_reg_60__1_ ( .D(n4438), .CLK(clk), .Q(arr[961]) );
  DFFPOSX1 arr_reg_60__0_ ( .D(n4437), .CLK(clk), .Q(arr[960]) );
  DFFPOSX1 arr_reg_59__15_ ( .D(n4436), .CLK(clk), .Q(arr[959]) );
  DFFPOSX1 arr_reg_59__14_ ( .D(n4435), .CLK(clk), .Q(arr[958]) );
  DFFPOSX1 arr_reg_59__13_ ( .D(n4434), .CLK(clk), .Q(arr[957]) );
  DFFPOSX1 arr_reg_59__12_ ( .D(n4433), .CLK(clk), .Q(arr[956]) );
  DFFPOSX1 arr_reg_59__11_ ( .D(n4432), .CLK(clk), .Q(arr[955]) );
  DFFPOSX1 arr_reg_59__10_ ( .D(n4431), .CLK(clk), .Q(arr[954]) );
  DFFPOSX1 arr_reg_59__9_ ( .D(n4430), .CLK(clk), .Q(arr[953]) );
  DFFPOSX1 arr_reg_59__8_ ( .D(n4429), .CLK(clk), .Q(arr[952]) );
  DFFPOSX1 arr_reg_59__7_ ( .D(n4428), .CLK(clk), .Q(arr[951]) );
  DFFPOSX1 arr_reg_59__6_ ( .D(n4427), .CLK(clk), .Q(arr[950]) );
  DFFPOSX1 arr_reg_59__5_ ( .D(n4426), .CLK(clk), .Q(arr[949]) );
  DFFPOSX1 arr_reg_59__4_ ( .D(n4425), .CLK(clk), .Q(arr[948]) );
  DFFPOSX1 arr_reg_59__3_ ( .D(n4424), .CLK(clk), .Q(arr[947]) );
  DFFPOSX1 arr_reg_59__2_ ( .D(n4423), .CLK(clk), .Q(arr[946]) );
  DFFPOSX1 arr_reg_59__1_ ( .D(n4422), .CLK(clk), .Q(arr[945]) );
  DFFPOSX1 arr_reg_59__0_ ( .D(n4421), .CLK(clk), .Q(arr[944]) );
  DFFPOSX1 arr_reg_58__15_ ( .D(n4420), .CLK(clk), .Q(arr[943]) );
  DFFPOSX1 arr_reg_58__14_ ( .D(n4419), .CLK(clk), .Q(arr[942]) );
  DFFPOSX1 arr_reg_58__13_ ( .D(n4418), .CLK(clk), .Q(arr[941]) );
  DFFPOSX1 arr_reg_58__12_ ( .D(n4417), .CLK(clk), .Q(arr[940]) );
  DFFPOSX1 arr_reg_58__11_ ( .D(n4416), .CLK(clk), .Q(arr[939]) );
  DFFPOSX1 arr_reg_58__10_ ( .D(n4415), .CLK(clk), .Q(arr[938]) );
  DFFPOSX1 arr_reg_58__9_ ( .D(n4414), .CLK(clk), .Q(arr[937]) );
  DFFPOSX1 arr_reg_58__8_ ( .D(n4413), .CLK(clk), .Q(arr[936]) );
  DFFPOSX1 arr_reg_58__7_ ( .D(n4412), .CLK(clk), .Q(arr[935]) );
  DFFPOSX1 arr_reg_58__6_ ( .D(n4411), .CLK(clk), .Q(arr[934]) );
  DFFPOSX1 arr_reg_58__5_ ( .D(n4410), .CLK(clk), .Q(arr[933]) );
  DFFPOSX1 arr_reg_58__4_ ( .D(n4409), .CLK(clk), .Q(arr[932]) );
  DFFPOSX1 arr_reg_58__3_ ( .D(n4408), .CLK(clk), .Q(arr[931]) );
  DFFPOSX1 arr_reg_58__2_ ( .D(n4407), .CLK(clk), .Q(arr[930]) );
  DFFPOSX1 arr_reg_58__1_ ( .D(n4406), .CLK(clk), .Q(arr[929]) );
  DFFPOSX1 arr_reg_58__0_ ( .D(n4405), .CLK(clk), .Q(arr[928]) );
  DFFPOSX1 arr_reg_57__15_ ( .D(n4404), .CLK(clk), .Q(arr[927]) );
  DFFPOSX1 arr_reg_57__14_ ( .D(n4403), .CLK(clk), .Q(arr[926]) );
  DFFPOSX1 arr_reg_57__13_ ( .D(n4402), .CLK(clk), .Q(arr[925]) );
  DFFPOSX1 arr_reg_57__12_ ( .D(n4401), .CLK(clk), .Q(arr[924]) );
  DFFPOSX1 arr_reg_57__11_ ( .D(n4400), .CLK(clk), .Q(arr[923]) );
  DFFPOSX1 arr_reg_57__10_ ( .D(n4399), .CLK(clk), .Q(arr[922]) );
  DFFPOSX1 arr_reg_57__9_ ( .D(n4398), .CLK(clk), .Q(arr[921]) );
  DFFPOSX1 arr_reg_57__8_ ( .D(n4397), .CLK(clk), .Q(arr[920]) );
  DFFPOSX1 arr_reg_57__7_ ( .D(n4396), .CLK(clk), .Q(arr[919]) );
  DFFPOSX1 arr_reg_57__6_ ( .D(n4395), .CLK(clk), .Q(arr[918]) );
  DFFPOSX1 arr_reg_57__5_ ( .D(n4394), .CLK(clk), .Q(arr[917]) );
  DFFPOSX1 arr_reg_57__4_ ( .D(n4393), .CLK(clk), .Q(arr[916]) );
  DFFPOSX1 arr_reg_57__3_ ( .D(n4392), .CLK(clk), .Q(arr[915]) );
  DFFPOSX1 arr_reg_57__2_ ( .D(n4391), .CLK(clk), .Q(arr[914]) );
  DFFPOSX1 arr_reg_57__1_ ( .D(n4390), .CLK(clk), .Q(arr[913]) );
  DFFPOSX1 arr_reg_57__0_ ( .D(n4389), .CLK(clk), .Q(arr[912]) );
  DFFPOSX1 arr_reg_56__15_ ( .D(n4388), .CLK(clk), .Q(arr[911]) );
  DFFPOSX1 arr_reg_56__14_ ( .D(n4387), .CLK(clk), .Q(arr[910]) );
  DFFPOSX1 arr_reg_56__13_ ( .D(n4386), .CLK(clk), .Q(arr[909]) );
  DFFPOSX1 arr_reg_56__12_ ( .D(n4385), .CLK(clk), .Q(arr[908]) );
  DFFPOSX1 arr_reg_56__11_ ( .D(n4384), .CLK(clk), .Q(arr[907]) );
  DFFPOSX1 arr_reg_56__10_ ( .D(n4383), .CLK(clk), .Q(arr[906]) );
  DFFPOSX1 arr_reg_56__9_ ( .D(n4382), .CLK(clk), .Q(arr[905]) );
  DFFPOSX1 arr_reg_56__8_ ( .D(n4381), .CLK(clk), .Q(arr[904]) );
  DFFPOSX1 arr_reg_56__7_ ( .D(n4380), .CLK(clk), .Q(arr[903]) );
  DFFPOSX1 arr_reg_56__6_ ( .D(n4379), .CLK(clk), .Q(arr[902]) );
  DFFPOSX1 arr_reg_56__5_ ( .D(n4378), .CLK(clk), .Q(arr[901]) );
  DFFPOSX1 arr_reg_56__4_ ( .D(n4377), .CLK(clk), .Q(arr[900]) );
  DFFPOSX1 arr_reg_56__3_ ( .D(n4376), .CLK(clk), .Q(arr[899]) );
  DFFPOSX1 arr_reg_56__2_ ( .D(n4375), .CLK(clk), .Q(arr[898]) );
  DFFPOSX1 arr_reg_56__1_ ( .D(n4374), .CLK(clk), .Q(arr[897]) );
  DFFPOSX1 arr_reg_56__0_ ( .D(n4373), .CLK(clk), .Q(arr[896]) );
  DFFPOSX1 arr_reg_55__15_ ( .D(n4372), .CLK(clk), .Q(arr[895]) );
  DFFPOSX1 arr_reg_55__14_ ( .D(n4371), .CLK(clk), .Q(arr[894]) );
  DFFPOSX1 arr_reg_55__13_ ( .D(n4370), .CLK(clk), .Q(arr[893]) );
  DFFPOSX1 arr_reg_55__12_ ( .D(n4369), .CLK(clk), .Q(arr[892]) );
  DFFPOSX1 arr_reg_55__11_ ( .D(n4368), .CLK(clk), .Q(arr[891]) );
  DFFPOSX1 arr_reg_55__10_ ( .D(n4367), .CLK(clk), .Q(arr[890]) );
  DFFPOSX1 arr_reg_55__9_ ( .D(n4366), .CLK(clk), .Q(arr[889]) );
  DFFPOSX1 arr_reg_55__8_ ( .D(n4365), .CLK(clk), .Q(arr[888]) );
  DFFPOSX1 arr_reg_55__7_ ( .D(n4364), .CLK(clk), .Q(arr[887]) );
  DFFPOSX1 arr_reg_55__6_ ( .D(n4363), .CLK(clk), .Q(arr[886]) );
  DFFPOSX1 arr_reg_55__5_ ( .D(n4362), .CLK(clk), .Q(arr[885]) );
  DFFPOSX1 arr_reg_55__4_ ( .D(n4361), .CLK(clk), .Q(arr[884]) );
  DFFPOSX1 arr_reg_55__3_ ( .D(n4360), .CLK(clk), .Q(arr[883]) );
  DFFPOSX1 arr_reg_55__2_ ( .D(n4359), .CLK(clk), .Q(arr[882]) );
  DFFPOSX1 arr_reg_55__1_ ( .D(n4358), .CLK(clk), .Q(arr[881]) );
  DFFPOSX1 arr_reg_55__0_ ( .D(n4357), .CLK(clk), .Q(arr[880]) );
  DFFPOSX1 arr_reg_54__15_ ( .D(n4356), .CLK(clk), .Q(arr[879]) );
  DFFPOSX1 arr_reg_54__14_ ( .D(n4355), .CLK(clk), .Q(arr[878]) );
  DFFPOSX1 arr_reg_54__13_ ( .D(n4354), .CLK(clk), .Q(arr[877]) );
  DFFPOSX1 arr_reg_54__12_ ( .D(n4353), .CLK(clk), .Q(arr[876]) );
  DFFPOSX1 arr_reg_54__11_ ( .D(n4352), .CLK(clk), .Q(arr[875]) );
  DFFPOSX1 arr_reg_54__10_ ( .D(n4351), .CLK(clk), .Q(arr[874]) );
  DFFPOSX1 arr_reg_54__9_ ( .D(n4350), .CLK(clk), .Q(arr[873]) );
  DFFPOSX1 arr_reg_54__8_ ( .D(n4349), .CLK(clk), .Q(arr[872]) );
  DFFPOSX1 arr_reg_54__7_ ( .D(n4348), .CLK(clk), .Q(arr[871]) );
  DFFPOSX1 arr_reg_54__6_ ( .D(n4347), .CLK(clk), .Q(arr[870]) );
  DFFPOSX1 arr_reg_54__5_ ( .D(n4346), .CLK(clk), .Q(arr[869]) );
  DFFPOSX1 arr_reg_54__4_ ( .D(n4345), .CLK(clk), .Q(arr[868]) );
  DFFPOSX1 arr_reg_54__3_ ( .D(n4344), .CLK(clk), .Q(arr[867]) );
  DFFPOSX1 arr_reg_54__2_ ( .D(n4343), .CLK(clk), .Q(arr[866]) );
  DFFPOSX1 arr_reg_54__1_ ( .D(n4342), .CLK(clk), .Q(arr[865]) );
  DFFPOSX1 arr_reg_54__0_ ( .D(n4341), .CLK(clk), .Q(arr[864]) );
  DFFPOSX1 arr_reg_53__15_ ( .D(n4340), .CLK(clk), .Q(arr[863]) );
  DFFPOSX1 arr_reg_53__14_ ( .D(n4339), .CLK(clk), .Q(arr[862]) );
  DFFPOSX1 arr_reg_53__13_ ( .D(n4338), .CLK(clk), .Q(arr[861]) );
  DFFPOSX1 arr_reg_53__12_ ( .D(n4337), .CLK(clk), .Q(arr[860]) );
  DFFPOSX1 arr_reg_53__11_ ( .D(n4336), .CLK(clk), .Q(arr[859]) );
  DFFPOSX1 arr_reg_53__10_ ( .D(n4335), .CLK(clk), .Q(arr[858]) );
  DFFPOSX1 arr_reg_53__9_ ( .D(n4334), .CLK(clk), .Q(arr[857]) );
  DFFPOSX1 arr_reg_53__8_ ( .D(n4333), .CLK(clk), .Q(arr[856]) );
  DFFPOSX1 arr_reg_53__7_ ( .D(n4332), .CLK(clk), .Q(arr[855]) );
  DFFPOSX1 arr_reg_53__6_ ( .D(n4331), .CLK(clk), .Q(arr[854]) );
  DFFPOSX1 arr_reg_53__5_ ( .D(n4330), .CLK(clk), .Q(arr[853]) );
  DFFPOSX1 arr_reg_53__4_ ( .D(n4329), .CLK(clk), .Q(arr[852]) );
  DFFPOSX1 arr_reg_53__3_ ( .D(n4328), .CLK(clk), .Q(arr[851]) );
  DFFPOSX1 arr_reg_53__2_ ( .D(n4327), .CLK(clk), .Q(arr[850]) );
  DFFPOSX1 arr_reg_53__1_ ( .D(n4326), .CLK(clk), .Q(arr[849]) );
  DFFPOSX1 arr_reg_53__0_ ( .D(n4325), .CLK(clk), .Q(arr[848]) );
  DFFPOSX1 arr_reg_52__15_ ( .D(n4324), .CLK(clk), .Q(arr[847]) );
  DFFPOSX1 arr_reg_52__14_ ( .D(n4323), .CLK(clk), .Q(arr[846]) );
  DFFPOSX1 arr_reg_52__13_ ( .D(n4322), .CLK(clk), .Q(arr[845]) );
  DFFPOSX1 arr_reg_52__12_ ( .D(n4321), .CLK(clk), .Q(arr[844]) );
  DFFPOSX1 arr_reg_52__11_ ( .D(n4320), .CLK(clk), .Q(arr[843]) );
  DFFPOSX1 arr_reg_52__10_ ( .D(n4319), .CLK(clk), .Q(arr[842]) );
  DFFPOSX1 arr_reg_52__9_ ( .D(n4318), .CLK(clk), .Q(arr[841]) );
  DFFPOSX1 arr_reg_52__8_ ( .D(n4317), .CLK(clk), .Q(arr[840]) );
  DFFPOSX1 arr_reg_52__7_ ( .D(n4316), .CLK(clk), .Q(arr[839]) );
  DFFPOSX1 arr_reg_52__6_ ( .D(n4315), .CLK(clk), .Q(arr[838]) );
  DFFPOSX1 arr_reg_52__5_ ( .D(n4314), .CLK(clk), .Q(arr[837]) );
  DFFPOSX1 arr_reg_52__4_ ( .D(n4313), .CLK(clk), .Q(arr[836]) );
  DFFPOSX1 arr_reg_52__3_ ( .D(n4312), .CLK(clk), .Q(arr[835]) );
  DFFPOSX1 arr_reg_52__2_ ( .D(n4311), .CLK(clk), .Q(arr[834]) );
  DFFPOSX1 arr_reg_52__1_ ( .D(n4310), .CLK(clk), .Q(arr[833]) );
  DFFPOSX1 arr_reg_52__0_ ( .D(n4309), .CLK(clk), .Q(arr[832]) );
  DFFPOSX1 arr_reg_51__15_ ( .D(n4308), .CLK(clk), .Q(arr[831]) );
  DFFPOSX1 arr_reg_51__14_ ( .D(n4307), .CLK(clk), .Q(arr[830]) );
  DFFPOSX1 arr_reg_51__13_ ( .D(n4306), .CLK(clk), .Q(arr[829]) );
  DFFPOSX1 arr_reg_51__12_ ( .D(n4305), .CLK(clk), .Q(arr[828]) );
  DFFPOSX1 arr_reg_51__11_ ( .D(n4304), .CLK(clk), .Q(arr[827]) );
  DFFPOSX1 arr_reg_51__10_ ( .D(n4303), .CLK(clk), .Q(arr[826]) );
  DFFPOSX1 arr_reg_51__9_ ( .D(n4302), .CLK(clk), .Q(arr[825]) );
  DFFPOSX1 arr_reg_51__8_ ( .D(n4301), .CLK(clk), .Q(arr[824]) );
  DFFPOSX1 arr_reg_51__7_ ( .D(n4300), .CLK(clk), .Q(arr[823]) );
  DFFPOSX1 arr_reg_51__6_ ( .D(n4299), .CLK(clk), .Q(arr[822]) );
  DFFPOSX1 arr_reg_51__5_ ( .D(n4298), .CLK(clk), .Q(arr[821]) );
  DFFPOSX1 arr_reg_51__4_ ( .D(n4297), .CLK(clk), .Q(arr[820]) );
  DFFPOSX1 arr_reg_51__3_ ( .D(n4296), .CLK(clk), .Q(arr[819]) );
  DFFPOSX1 arr_reg_51__2_ ( .D(n4295), .CLK(clk), .Q(arr[818]) );
  DFFPOSX1 arr_reg_51__1_ ( .D(n4294), .CLK(clk), .Q(arr[817]) );
  DFFPOSX1 arr_reg_51__0_ ( .D(n4293), .CLK(clk), .Q(arr[816]) );
  DFFPOSX1 arr_reg_50__15_ ( .D(n4292), .CLK(clk), .Q(arr[815]) );
  DFFPOSX1 arr_reg_50__14_ ( .D(n4291), .CLK(clk), .Q(arr[814]) );
  DFFPOSX1 arr_reg_50__13_ ( .D(n4290), .CLK(clk), .Q(arr[813]) );
  DFFPOSX1 arr_reg_50__12_ ( .D(n4289), .CLK(clk), .Q(arr[812]) );
  DFFPOSX1 arr_reg_50__11_ ( .D(n4288), .CLK(clk), .Q(arr[811]) );
  DFFPOSX1 arr_reg_50__10_ ( .D(n4287), .CLK(clk), .Q(arr[810]) );
  DFFPOSX1 arr_reg_50__9_ ( .D(n4286), .CLK(clk), .Q(arr[809]) );
  DFFPOSX1 arr_reg_50__8_ ( .D(n4285), .CLK(clk), .Q(arr[808]) );
  DFFPOSX1 arr_reg_50__7_ ( .D(n4284), .CLK(clk), .Q(arr[807]) );
  DFFPOSX1 arr_reg_50__6_ ( .D(n4283), .CLK(clk), .Q(arr[806]) );
  DFFPOSX1 arr_reg_50__5_ ( .D(n4282), .CLK(clk), .Q(arr[805]) );
  DFFPOSX1 arr_reg_50__4_ ( .D(n4281), .CLK(clk), .Q(arr[804]) );
  DFFPOSX1 arr_reg_50__3_ ( .D(n4280), .CLK(clk), .Q(arr[803]) );
  DFFPOSX1 arr_reg_50__2_ ( .D(n4279), .CLK(clk), .Q(arr[802]) );
  DFFPOSX1 arr_reg_50__1_ ( .D(n4278), .CLK(clk), .Q(arr[801]) );
  DFFPOSX1 arr_reg_50__0_ ( .D(n4277), .CLK(clk), .Q(arr[800]) );
  DFFPOSX1 arr_reg_49__15_ ( .D(n4276), .CLK(clk), .Q(arr[799]) );
  DFFPOSX1 arr_reg_49__14_ ( .D(n4275), .CLK(clk), .Q(arr[798]) );
  DFFPOSX1 arr_reg_49__13_ ( .D(n4274), .CLK(clk), .Q(arr[797]) );
  DFFPOSX1 arr_reg_49__12_ ( .D(n4273), .CLK(clk), .Q(arr[796]) );
  DFFPOSX1 arr_reg_49__11_ ( .D(n4272), .CLK(clk), .Q(arr[795]) );
  DFFPOSX1 arr_reg_49__10_ ( .D(n4271), .CLK(clk), .Q(arr[794]) );
  DFFPOSX1 arr_reg_49__9_ ( .D(n4270), .CLK(clk), .Q(arr[793]) );
  DFFPOSX1 arr_reg_49__8_ ( .D(n4269), .CLK(clk), .Q(arr[792]) );
  DFFPOSX1 arr_reg_49__7_ ( .D(n4268), .CLK(clk), .Q(arr[791]) );
  DFFPOSX1 arr_reg_49__6_ ( .D(n4267), .CLK(clk), .Q(arr[790]) );
  DFFPOSX1 arr_reg_49__5_ ( .D(n4266), .CLK(clk), .Q(arr[789]) );
  DFFPOSX1 arr_reg_49__4_ ( .D(n4265), .CLK(clk), .Q(arr[788]) );
  DFFPOSX1 arr_reg_49__3_ ( .D(n4264), .CLK(clk), .Q(arr[787]) );
  DFFPOSX1 arr_reg_49__2_ ( .D(n4263), .CLK(clk), .Q(arr[786]) );
  DFFPOSX1 arr_reg_49__1_ ( .D(n4262), .CLK(clk), .Q(arr[785]) );
  DFFPOSX1 arr_reg_49__0_ ( .D(n4261), .CLK(clk), .Q(arr[784]) );
  DFFPOSX1 arr_reg_48__15_ ( .D(n4260), .CLK(clk), .Q(arr[783]) );
  DFFPOSX1 arr_reg_48__14_ ( .D(n4259), .CLK(clk), .Q(arr[782]) );
  DFFPOSX1 arr_reg_48__13_ ( .D(n4258), .CLK(clk), .Q(arr[781]) );
  DFFPOSX1 arr_reg_48__12_ ( .D(n4257), .CLK(clk), .Q(arr[780]) );
  DFFPOSX1 arr_reg_48__11_ ( .D(n4256), .CLK(clk), .Q(arr[779]) );
  DFFPOSX1 arr_reg_48__10_ ( .D(n4255), .CLK(clk), .Q(arr[778]) );
  DFFPOSX1 arr_reg_48__9_ ( .D(n4254), .CLK(clk), .Q(arr[777]) );
  DFFPOSX1 arr_reg_48__8_ ( .D(n4253), .CLK(clk), .Q(arr[776]) );
  DFFPOSX1 arr_reg_48__7_ ( .D(n4252), .CLK(clk), .Q(arr[775]) );
  DFFPOSX1 arr_reg_48__6_ ( .D(n4251), .CLK(clk), .Q(arr[774]) );
  DFFPOSX1 arr_reg_48__5_ ( .D(n4250), .CLK(clk), .Q(arr[773]) );
  DFFPOSX1 arr_reg_48__4_ ( .D(n4249), .CLK(clk), .Q(arr[772]) );
  DFFPOSX1 arr_reg_48__3_ ( .D(n4248), .CLK(clk), .Q(arr[771]) );
  DFFPOSX1 arr_reg_48__2_ ( .D(n4247), .CLK(clk), .Q(arr[770]) );
  DFFPOSX1 arr_reg_48__1_ ( .D(n4246), .CLK(clk), .Q(arr[769]) );
  DFFPOSX1 arr_reg_48__0_ ( .D(n4245), .CLK(clk), .Q(arr[768]) );
  DFFPOSX1 arr_reg_47__15_ ( .D(n4244), .CLK(clk), .Q(arr[767]) );
  DFFPOSX1 arr_reg_47__14_ ( .D(n4243), .CLK(clk), .Q(arr[766]) );
  DFFPOSX1 arr_reg_47__13_ ( .D(n4242), .CLK(clk), .Q(arr[765]) );
  DFFPOSX1 arr_reg_47__12_ ( .D(n4241), .CLK(clk), .Q(arr[764]) );
  DFFPOSX1 arr_reg_47__11_ ( .D(n4240), .CLK(clk), .Q(arr[763]) );
  DFFPOSX1 arr_reg_47__10_ ( .D(n4239), .CLK(clk), .Q(arr[762]) );
  DFFPOSX1 arr_reg_47__9_ ( .D(n4238), .CLK(clk), .Q(arr[761]) );
  DFFPOSX1 arr_reg_47__8_ ( .D(n4237), .CLK(clk), .Q(arr[760]) );
  DFFPOSX1 arr_reg_47__7_ ( .D(n4236), .CLK(clk), .Q(arr[759]) );
  DFFPOSX1 arr_reg_47__6_ ( .D(n4235), .CLK(clk), .Q(arr[758]) );
  DFFPOSX1 arr_reg_47__5_ ( .D(n4234), .CLK(clk), .Q(arr[757]) );
  DFFPOSX1 arr_reg_47__4_ ( .D(n4233), .CLK(clk), .Q(arr[756]) );
  DFFPOSX1 arr_reg_47__3_ ( .D(n4232), .CLK(clk), .Q(arr[755]) );
  DFFPOSX1 arr_reg_47__2_ ( .D(n4231), .CLK(clk), .Q(arr[754]) );
  DFFPOSX1 arr_reg_47__1_ ( .D(n4230), .CLK(clk), .Q(arr[753]) );
  DFFPOSX1 arr_reg_47__0_ ( .D(n4229), .CLK(clk), .Q(arr[752]) );
  DFFPOSX1 arr_reg_46__15_ ( .D(n4228), .CLK(clk), .Q(arr[751]) );
  DFFPOSX1 arr_reg_46__14_ ( .D(n4227), .CLK(clk), .Q(arr[750]) );
  DFFPOSX1 arr_reg_46__13_ ( .D(n4226), .CLK(clk), .Q(arr[749]) );
  DFFPOSX1 arr_reg_46__12_ ( .D(n4225), .CLK(clk), .Q(arr[748]) );
  DFFPOSX1 arr_reg_46__11_ ( .D(n4224), .CLK(clk), .Q(arr[747]) );
  DFFPOSX1 arr_reg_46__10_ ( .D(n4223), .CLK(clk), .Q(arr[746]) );
  DFFPOSX1 arr_reg_46__9_ ( .D(n4222), .CLK(clk), .Q(arr[745]) );
  DFFPOSX1 arr_reg_46__8_ ( .D(n4221), .CLK(clk), .Q(arr[744]) );
  DFFPOSX1 arr_reg_46__7_ ( .D(n4220), .CLK(clk), .Q(arr[743]) );
  DFFPOSX1 arr_reg_46__6_ ( .D(n4219), .CLK(clk), .Q(arr[742]) );
  DFFPOSX1 arr_reg_46__5_ ( .D(n4218), .CLK(clk), .Q(arr[741]) );
  DFFPOSX1 arr_reg_46__4_ ( .D(n4217), .CLK(clk), .Q(arr[740]) );
  DFFPOSX1 arr_reg_46__3_ ( .D(n4216), .CLK(clk), .Q(arr[739]) );
  DFFPOSX1 arr_reg_46__2_ ( .D(n4215), .CLK(clk), .Q(arr[738]) );
  DFFPOSX1 arr_reg_46__1_ ( .D(n4214), .CLK(clk), .Q(arr[737]) );
  DFFPOSX1 arr_reg_46__0_ ( .D(n4213), .CLK(clk), .Q(arr[736]) );
  DFFPOSX1 arr_reg_45__15_ ( .D(n4212), .CLK(clk), .Q(arr[735]) );
  DFFPOSX1 arr_reg_45__14_ ( .D(n4211), .CLK(clk), .Q(arr[734]) );
  DFFPOSX1 arr_reg_45__13_ ( .D(n4210), .CLK(clk), .Q(arr[733]) );
  DFFPOSX1 arr_reg_45__12_ ( .D(n4209), .CLK(clk), .Q(arr[732]) );
  DFFPOSX1 arr_reg_45__11_ ( .D(n4208), .CLK(clk), .Q(arr[731]) );
  DFFPOSX1 arr_reg_45__10_ ( .D(n4207), .CLK(clk), .Q(arr[730]) );
  DFFPOSX1 arr_reg_45__9_ ( .D(n4206), .CLK(clk), .Q(arr[729]) );
  DFFPOSX1 arr_reg_45__8_ ( .D(n4205), .CLK(clk), .Q(arr[728]) );
  DFFPOSX1 arr_reg_45__7_ ( .D(n4204), .CLK(clk), .Q(arr[727]) );
  DFFPOSX1 arr_reg_45__6_ ( .D(n4203), .CLK(clk), .Q(arr[726]) );
  DFFPOSX1 arr_reg_45__5_ ( .D(n4202), .CLK(clk), .Q(arr[725]) );
  DFFPOSX1 arr_reg_45__4_ ( .D(n4201), .CLK(clk), .Q(arr[724]) );
  DFFPOSX1 arr_reg_45__3_ ( .D(n4200), .CLK(clk), .Q(arr[723]) );
  DFFPOSX1 arr_reg_45__2_ ( .D(n4199), .CLK(clk), .Q(arr[722]) );
  DFFPOSX1 arr_reg_45__1_ ( .D(n4198), .CLK(clk), .Q(arr[721]) );
  DFFPOSX1 arr_reg_45__0_ ( .D(n4197), .CLK(clk), .Q(arr[720]) );
  DFFPOSX1 arr_reg_44__15_ ( .D(n4196), .CLK(clk), .Q(arr[719]) );
  DFFPOSX1 arr_reg_44__14_ ( .D(n4195), .CLK(clk), .Q(arr[718]) );
  DFFPOSX1 arr_reg_44__13_ ( .D(n4194), .CLK(clk), .Q(arr[717]) );
  DFFPOSX1 arr_reg_44__12_ ( .D(n4193), .CLK(clk), .Q(arr[716]) );
  DFFPOSX1 arr_reg_44__11_ ( .D(n4192), .CLK(clk), .Q(arr[715]) );
  DFFPOSX1 arr_reg_44__10_ ( .D(n4191), .CLK(clk), .Q(arr[714]) );
  DFFPOSX1 arr_reg_44__9_ ( .D(n4190), .CLK(clk), .Q(arr[713]) );
  DFFPOSX1 arr_reg_44__8_ ( .D(n4189), .CLK(clk), .Q(arr[712]) );
  DFFPOSX1 arr_reg_44__7_ ( .D(n4188), .CLK(clk), .Q(arr[711]) );
  DFFPOSX1 arr_reg_44__6_ ( .D(n4187), .CLK(clk), .Q(arr[710]) );
  DFFPOSX1 arr_reg_44__5_ ( .D(n4186), .CLK(clk), .Q(arr[709]) );
  DFFPOSX1 arr_reg_44__4_ ( .D(n4185), .CLK(clk), .Q(arr[708]) );
  DFFPOSX1 arr_reg_44__3_ ( .D(n4184), .CLK(clk), .Q(arr[707]) );
  DFFPOSX1 arr_reg_44__2_ ( .D(n4183), .CLK(clk), .Q(arr[706]) );
  DFFPOSX1 arr_reg_44__1_ ( .D(n4182), .CLK(clk), .Q(arr[705]) );
  DFFPOSX1 arr_reg_44__0_ ( .D(n4181), .CLK(clk), .Q(arr[704]) );
  DFFPOSX1 arr_reg_43__15_ ( .D(n4180), .CLK(clk), .Q(arr[703]) );
  DFFPOSX1 arr_reg_43__14_ ( .D(n4179), .CLK(clk), .Q(arr[702]) );
  DFFPOSX1 arr_reg_43__13_ ( .D(n4178), .CLK(clk), .Q(arr[701]) );
  DFFPOSX1 arr_reg_43__12_ ( .D(n4177), .CLK(clk), .Q(arr[700]) );
  DFFPOSX1 arr_reg_43__11_ ( .D(n4176), .CLK(clk), .Q(arr[699]) );
  DFFPOSX1 arr_reg_43__10_ ( .D(n4175), .CLK(clk), .Q(arr[698]) );
  DFFPOSX1 arr_reg_43__9_ ( .D(n4174), .CLK(clk), .Q(arr[697]) );
  DFFPOSX1 arr_reg_43__8_ ( .D(n4173), .CLK(clk), .Q(arr[696]) );
  DFFPOSX1 arr_reg_43__7_ ( .D(n4172), .CLK(clk), .Q(arr[695]) );
  DFFPOSX1 arr_reg_43__6_ ( .D(n4171), .CLK(clk), .Q(arr[694]) );
  DFFPOSX1 arr_reg_43__5_ ( .D(n4170), .CLK(clk), .Q(arr[693]) );
  DFFPOSX1 arr_reg_43__4_ ( .D(n4169), .CLK(clk), .Q(arr[692]) );
  DFFPOSX1 arr_reg_43__3_ ( .D(n4168), .CLK(clk), .Q(arr[691]) );
  DFFPOSX1 arr_reg_43__2_ ( .D(n4167), .CLK(clk), .Q(arr[690]) );
  DFFPOSX1 arr_reg_43__1_ ( .D(n4166), .CLK(clk), .Q(arr[689]) );
  DFFPOSX1 arr_reg_43__0_ ( .D(n4165), .CLK(clk), .Q(arr[688]) );
  DFFPOSX1 arr_reg_42__15_ ( .D(n4164), .CLK(clk), .Q(arr[687]) );
  DFFPOSX1 arr_reg_42__14_ ( .D(n4163), .CLK(clk), .Q(arr[686]) );
  DFFPOSX1 arr_reg_42__13_ ( .D(n4162), .CLK(clk), .Q(arr[685]) );
  DFFPOSX1 arr_reg_42__12_ ( .D(n4161), .CLK(clk), .Q(arr[684]) );
  DFFPOSX1 arr_reg_42__11_ ( .D(n4160), .CLK(clk), .Q(arr[683]) );
  DFFPOSX1 arr_reg_42__10_ ( .D(n4159), .CLK(clk), .Q(arr[682]) );
  DFFPOSX1 arr_reg_42__9_ ( .D(n4158), .CLK(clk), .Q(arr[681]) );
  DFFPOSX1 arr_reg_42__8_ ( .D(n4157), .CLK(clk), .Q(arr[680]) );
  DFFPOSX1 arr_reg_42__7_ ( .D(n4156), .CLK(clk), .Q(arr[679]) );
  DFFPOSX1 arr_reg_42__6_ ( .D(n4155), .CLK(clk), .Q(arr[678]) );
  DFFPOSX1 arr_reg_42__5_ ( .D(n4154), .CLK(clk), .Q(arr[677]) );
  DFFPOSX1 arr_reg_42__4_ ( .D(n4153), .CLK(clk), .Q(arr[676]) );
  DFFPOSX1 arr_reg_42__3_ ( .D(n4152), .CLK(clk), .Q(arr[675]) );
  DFFPOSX1 arr_reg_42__2_ ( .D(n4151), .CLK(clk), .Q(arr[674]) );
  DFFPOSX1 arr_reg_42__1_ ( .D(n4150), .CLK(clk), .Q(arr[673]) );
  DFFPOSX1 arr_reg_42__0_ ( .D(n4149), .CLK(clk), .Q(arr[672]) );
  DFFPOSX1 arr_reg_41__15_ ( .D(n4148), .CLK(clk), .Q(arr[671]) );
  DFFPOSX1 arr_reg_41__14_ ( .D(n4147), .CLK(clk), .Q(arr[670]) );
  DFFPOSX1 arr_reg_41__13_ ( .D(n4146), .CLK(clk), .Q(arr[669]) );
  DFFPOSX1 arr_reg_41__12_ ( .D(n4145), .CLK(clk), .Q(arr[668]) );
  DFFPOSX1 arr_reg_41__11_ ( .D(n4144), .CLK(clk), .Q(arr[667]) );
  DFFPOSX1 arr_reg_41__10_ ( .D(n4143), .CLK(clk), .Q(arr[666]) );
  DFFPOSX1 arr_reg_41__9_ ( .D(n4142), .CLK(clk), .Q(arr[665]) );
  DFFPOSX1 arr_reg_41__8_ ( .D(n4141), .CLK(clk), .Q(arr[664]) );
  DFFPOSX1 arr_reg_41__7_ ( .D(n4140), .CLK(clk), .Q(arr[663]) );
  DFFPOSX1 arr_reg_41__6_ ( .D(n4139), .CLK(clk), .Q(arr[662]) );
  DFFPOSX1 arr_reg_41__5_ ( .D(n4138), .CLK(clk), .Q(arr[661]) );
  DFFPOSX1 arr_reg_41__4_ ( .D(n4137), .CLK(clk), .Q(arr[660]) );
  DFFPOSX1 arr_reg_41__3_ ( .D(n4136), .CLK(clk), .Q(arr[659]) );
  DFFPOSX1 arr_reg_41__2_ ( .D(n4135), .CLK(clk), .Q(arr[658]) );
  DFFPOSX1 arr_reg_41__1_ ( .D(n4134), .CLK(clk), .Q(arr[657]) );
  DFFPOSX1 arr_reg_41__0_ ( .D(n4133), .CLK(clk), .Q(arr[656]) );
  DFFPOSX1 arr_reg_40__15_ ( .D(n4132), .CLK(clk), .Q(arr[655]) );
  DFFPOSX1 arr_reg_40__14_ ( .D(n4131), .CLK(clk), .Q(arr[654]) );
  DFFPOSX1 arr_reg_40__13_ ( .D(n4130), .CLK(clk), .Q(arr[653]) );
  DFFPOSX1 arr_reg_40__12_ ( .D(n4129), .CLK(clk), .Q(arr[652]) );
  DFFPOSX1 arr_reg_40__11_ ( .D(n4128), .CLK(clk), .Q(arr[651]) );
  DFFPOSX1 arr_reg_40__10_ ( .D(n4127), .CLK(clk), .Q(arr[650]) );
  DFFPOSX1 arr_reg_40__9_ ( .D(n4126), .CLK(clk), .Q(arr[649]) );
  DFFPOSX1 arr_reg_40__8_ ( .D(n4125), .CLK(clk), .Q(arr[648]) );
  DFFPOSX1 arr_reg_40__7_ ( .D(n4124), .CLK(clk), .Q(arr[647]) );
  DFFPOSX1 arr_reg_40__6_ ( .D(n4123), .CLK(clk), .Q(arr[646]) );
  DFFPOSX1 arr_reg_40__5_ ( .D(n4122), .CLK(clk), .Q(arr[645]) );
  DFFPOSX1 arr_reg_40__4_ ( .D(n4121), .CLK(clk), .Q(arr[644]) );
  DFFPOSX1 arr_reg_40__3_ ( .D(n4120), .CLK(clk), .Q(arr[643]) );
  DFFPOSX1 arr_reg_40__2_ ( .D(n4119), .CLK(clk), .Q(arr[642]) );
  DFFPOSX1 arr_reg_40__1_ ( .D(n4118), .CLK(clk), .Q(arr[641]) );
  DFFPOSX1 arr_reg_40__0_ ( .D(n4117), .CLK(clk), .Q(arr[640]) );
  DFFPOSX1 arr_reg_39__15_ ( .D(n4116), .CLK(clk), .Q(arr[639]) );
  DFFPOSX1 arr_reg_39__14_ ( .D(n4115), .CLK(clk), .Q(arr[638]) );
  DFFPOSX1 arr_reg_39__13_ ( .D(n4114), .CLK(clk), .Q(arr[637]) );
  DFFPOSX1 arr_reg_39__12_ ( .D(n4113), .CLK(clk), .Q(arr[636]) );
  DFFPOSX1 arr_reg_39__11_ ( .D(n4112), .CLK(clk), .Q(arr[635]) );
  DFFPOSX1 arr_reg_39__10_ ( .D(n4111), .CLK(clk), .Q(arr[634]) );
  DFFPOSX1 arr_reg_39__9_ ( .D(n4110), .CLK(clk), .Q(arr[633]) );
  DFFPOSX1 arr_reg_39__8_ ( .D(n4109), .CLK(clk), .Q(arr[632]) );
  DFFPOSX1 arr_reg_39__7_ ( .D(n4108), .CLK(clk), .Q(arr[631]) );
  DFFPOSX1 arr_reg_39__6_ ( .D(n4107), .CLK(clk), .Q(arr[630]) );
  DFFPOSX1 arr_reg_39__5_ ( .D(n4106), .CLK(clk), .Q(arr[629]) );
  DFFPOSX1 arr_reg_39__4_ ( .D(n4105), .CLK(clk), .Q(arr[628]) );
  DFFPOSX1 arr_reg_39__3_ ( .D(n4104), .CLK(clk), .Q(arr[627]) );
  DFFPOSX1 arr_reg_39__2_ ( .D(n4103), .CLK(clk), .Q(arr[626]) );
  DFFPOSX1 arr_reg_39__1_ ( .D(n4102), .CLK(clk), .Q(arr[625]) );
  DFFPOSX1 arr_reg_39__0_ ( .D(n4101), .CLK(clk), .Q(arr[624]) );
  DFFPOSX1 arr_reg_38__15_ ( .D(n4100), .CLK(clk), .Q(arr[623]) );
  DFFPOSX1 arr_reg_38__14_ ( .D(n4099), .CLK(clk), .Q(arr[622]) );
  DFFPOSX1 arr_reg_38__13_ ( .D(n4098), .CLK(clk), .Q(arr[621]) );
  DFFPOSX1 arr_reg_38__12_ ( .D(n4097), .CLK(clk), .Q(arr[620]) );
  DFFPOSX1 arr_reg_38__11_ ( .D(n4096), .CLK(clk), .Q(arr[619]) );
  DFFPOSX1 arr_reg_38__10_ ( .D(n4095), .CLK(clk), .Q(arr[618]) );
  DFFPOSX1 arr_reg_38__9_ ( .D(n4094), .CLK(clk), .Q(arr[617]) );
  DFFPOSX1 arr_reg_38__8_ ( .D(n4093), .CLK(clk), .Q(arr[616]) );
  DFFPOSX1 arr_reg_38__7_ ( .D(n4092), .CLK(clk), .Q(arr[615]) );
  DFFPOSX1 arr_reg_38__6_ ( .D(n4091), .CLK(clk), .Q(arr[614]) );
  DFFPOSX1 arr_reg_38__5_ ( .D(n4090), .CLK(clk), .Q(arr[613]) );
  DFFPOSX1 arr_reg_38__4_ ( .D(n4089), .CLK(clk), .Q(arr[612]) );
  DFFPOSX1 arr_reg_38__3_ ( .D(n4088), .CLK(clk), .Q(arr[611]) );
  DFFPOSX1 arr_reg_38__2_ ( .D(n4087), .CLK(clk), .Q(arr[610]) );
  DFFPOSX1 arr_reg_38__1_ ( .D(n4086), .CLK(clk), .Q(arr[609]) );
  DFFPOSX1 arr_reg_38__0_ ( .D(n4085), .CLK(clk), .Q(arr[608]) );
  DFFPOSX1 arr_reg_37__15_ ( .D(n4084), .CLK(clk), .Q(arr[607]) );
  DFFPOSX1 arr_reg_37__14_ ( .D(n4083), .CLK(clk), .Q(arr[606]) );
  DFFPOSX1 arr_reg_37__13_ ( .D(n4082), .CLK(clk), .Q(arr[605]) );
  DFFPOSX1 arr_reg_37__12_ ( .D(n4081), .CLK(clk), .Q(arr[604]) );
  DFFPOSX1 arr_reg_37__11_ ( .D(n4080), .CLK(clk), .Q(arr[603]) );
  DFFPOSX1 arr_reg_37__10_ ( .D(n4079), .CLK(clk), .Q(arr[602]) );
  DFFPOSX1 arr_reg_37__9_ ( .D(n4078), .CLK(clk), .Q(arr[601]) );
  DFFPOSX1 arr_reg_37__8_ ( .D(n4077), .CLK(clk), .Q(arr[600]) );
  DFFPOSX1 arr_reg_37__7_ ( .D(n4076), .CLK(clk), .Q(arr[599]) );
  DFFPOSX1 arr_reg_37__6_ ( .D(n4075), .CLK(clk), .Q(arr[598]) );
  DFFPOSX1 arr_reg_37__5_ ( .D(n4074), .CLK(clk), .Q(arr[597]) );
  DFFPOSX1 arr_reg_37__4_ ( .D(n4073), .CLK(clk), .Q(arr[596]) );
  DFFPOSX1 arr_reg_37__3_ ( .D(n4072), .CLK(clk), .Q(arr[595]) );
  DFFPOSX1 arr_reg_37__2_ ( .D(n4071), .CLK(clk), .Q(arr[594]) );
  DFFPOSX1 arr_reg_37__1_ ( .D(n4070), .CLK(clk), .Q(arr[593]) );
  DFFPOSX1 arr_reg_37__0_ ( .D(n4069), .CLK(clk), .Q(arr[592]) );
  DFFPOSX1 arr_reg_36__15_ ( .D(n4068), .CLK(clk), .Q(arr[591]) );
  DFFPOSX1 arr_reg_36__14_ ( .D(n4067), .CLK(clk), .Q(arr[590]) );
  DFFPOSX1 arr_reg_36__13_ ( .D(n4066), .CLK(clk), .Q(arr[589]) );
  DFFPOSX1 arr_reg_36__12_ ( .D(n4065), .CLK(clk), .Q(arr[588]) );
  DFFPOSX1 arr_reg_36__11_ ( .D(n4064), .CLK(clk), .Q(arr[587]) );
  DFFPOSX1 arr_reg_36__10_ ( .D(n4063), .CLK(clk), .Q(arr[586]) );
  DFFPOSX1 arr_reg_36__9_ ( .D(n4062), .CLK(clk), .Q(arr[585]) );
  DFFPOSX1 arr_reg_36__8_ ( .D(n4061), .CLK(clk), .Q(arr[584]) );
  DFFPOSX1 arr_reg_36__7_ ( .D(n4060), .CLK(clk), .Q(arr[583]) );
  DFFPOSX1 arr_reg_36__6_ ( .D(n4059), .CLK(clk), .Q(arr[582]) );
  DFFPOSX1 arr_reg_36__5_ ( .D(n4058), .CLK(clk), .Q(arr[581]) );
  DFFPOSX1 arr_reg_36__4_ ( .D(n4057), .CLK(clk), .Q(arr[580]) );
  DFFPOSX1 arr_reg_36__3_ ( .D(n4056), .CLK(clk), .Q(arr[579]) );
  DFFPOSX1 arr_reg_36__2_ ( .D(n4055), .CLK(clk), .Q(arr[578]) );
  DFFPOSX1 arr_reg_36__1_ ( .D(n4054), .CLK(clk), .Q(arr[577]) );
  DFFPOSX1 arr_reg_36__0_ ( .D(n4053), .CLK(clk), .Q(arr[576]) );
  DFFPOSX1 arr_reg_35__15_ ( .D(n4052), .CLK(clk), .Q(arr[575]) );
  DFFPOSX1 arr_reg_35__14_ ( .D(n4051), .CLK(clk), .Q(arr[574]) );
  DFFPOSX1 arr_reg_35__13_ ( .D(n4050), .CLK(clk), .Q(arr[573]) );
  DFFPOSX1 arr_reg_35__12_ ( .D(n4049), .CLK(clk), .Q(arr[572]) );
  DFFPOSX1 arr_reg_35__11_ ( .D(n4048), .CLK(clk), .Q(arr[571]) );
  DFFPOSX1 arr_reg_35__10_ ( .D(n4047), .CLK(clk), .Q(arr[570]) );
  DFFPOSX1 arr_reg_35__9_ ( .D(n4046), .CLK(clk), .Q(arr[569]) );
  DFFPOSX1 arr_reg_35__8_ ( .D(n4045), .CLK(clk), .Q(arr[568]) );
  DFFPOSX1 arr_reg_35__7_ ( .D(n4044), .CLK(clk), .Q(arr[567]) );
  DFFPOSX1 arr_reg_35__6_ ( .D(n4043), .CLK(clk), .Q(arr[566]) );
  DFFPOSX1 arr_reg_35__5_ ( .D(n4042), .CLK(clk), .Q(arr[565]) );
  DFFPOSX1 arr_reg_35__4_ ( .D(n4041), .CLK(clk), .Q(arr[564]) );
  DFFPOSX1 arr_reg_35__3_ ( .D(n4040), .CLK(clk), .Q(arr[563]) );
  DFFPOSX1 arr_reg_35__2_ ( .D(n4039), .CLK(clk), .Q(arr[562]) );
  DFFPOSX1 arr_reg_35__1_ ( .D(n4038), .CLK(clk), .Q(arr[561]) );
  DFFPOSX1 arr_reg_35__0_ ( .D(n4037), .CLK(clk), .Q(arr[560]) );
  DFFPOSX1 arr_reg_34__15_ ( .D(n4036), .CLK(clk), .Q(arr[559]) );
  DFFPOSX1 arr_reg_34__14_ ( .D(n4035), .CLK(clk), .Q(arr[558]) );
  DFFPOSX1 arr_reg_34__13_ ( .D(n4034), .CLK(clk), .Q(arr[557]) );
  DFFPOSX1 arr_reg_34__12_ ( .D(n4033), .CLK(clk), .Q(arr[556]) );
  DFFPOSX1 arr_reg_34__11_ ( .D(n4032), .CLK(clk), .Q(arr[555]) );
  DFFPOSX1 arr_reg_34__10_ ( .D(n4031), .CLK(clk), .Q(arr[554]) );
  DFFPOSX1 arr_reg_34__9_ ( .D(n4030), .CLK(clk), .Q(arr[553]) );
  DFFPOSX1 arr_reg_34__8_ ( .D(n4029), .CLK(clk), .Q(arr[552]) );
  DFFPOSX1 arr_reg_34__7_ ( .D(n4028), .CLK(clk), .Q(arr[551]) );
  DFFPOSX1 arr_reg_34__6_ ( .D(n4027), .CLK(clk), .Q(arr[550]) );
  DFFPOSX1 arr_reg_34__5_ ( .D(n4026), .CLK(clk), .Q(arr[549]) );
  DFFPOSX1 arr_reg_34__4_ ( .D(n4025), .CLK(clk), .Q(arr[548]) );
  DFFPOSX1 arr_reg_34__3_ ( .D(n4024), .CLK(clk), .Q(arr[547]) );
  DFFPOSX1 arr_reg_34__2_ ( .D(n4023), .CLK(clk), .Q(arr[546]) );
  DFFPOSX1 arr_reg_34__1_ ( .D(n4022), .CLK(clk), .Q(arr[545]) );
  DFFPOSX1 arr_reg_34__0_ ( .D(n4021), .CLK(clk), .Q(arr[544]) );
  DFFPOSX1 arr_reg_33__15_ ( .D(n4020), .CLK(clk), .Q(arr[543]) );
  DFFPOSX1 arr_reg_33__14_ ( .D(n4019), .CLK(clk), .Q(arr[542]) );
  DFFPOSX1 arr_reg_33__13_ ( .D(n4018), .CLK(clk), .Q(arr[541]) );
  DFFPOSX1 arr_reg_33__12_ ( .D(n4017), .CLK(clk), .Q(arr[540]) );
  DFFPOSX1 arr_reg_33__11_ ( .D(n4016), .CLK(clk), .Q(arr[539]) );
  DFFPOSX1 arr_reg_33__10_ ( .D(n4015), .CLK(clk), .Q(arr[538]) );
  DFFPOSX1 arr_reg_33__9_ ( .D(n4014), .CLK(clk), .Q(arr[537]) );
  DFFPOSX1 arr_reg_33__8_ ( .D(n4013), .CLK(clk), .Q(arr[536]) );
  DFFPOSX1 arr_reg_33__7_ ( .D(n4012), .CLK(clk), .Q(arr[535]) );
  DFFPOSX1 arr_reg_33__6_ ( .D(n4011), .CLK(clk), .Q(arr[534]) );
  DFFPOSX1 arr_reg_33__5_ ( .D(n4010), .CLK(clk), .Q(arr[533]) );
  DFFPOSX1 arr_reg_33__4_ ( .D(n4009), .CLK(clk), .Q(arr[532]) );
  DFFPOSX1 arr_reg_33__3_ ( .D(n4008), .CLK(clk), .Q(arr[531]) );
  DFFPOSX1 arr_reg_33__2_ ( .D(n4007), .CLK(clk), .Q(arr[530]) );
  DFFPOSX1 arr_reg_33__1_ ( .D(n4006), .CLK(clk), .Q(arr[529]) );
  DFFPOSX1 arr_reg_33__0_ ( .D(n4005), .CLK(clk), .Q(arr[528]) );
  DFFPOSX1 arr_reg_32__15_ ( .D(n4004), .CLK(clk), .Q(arr[527]) );
  DFFPOSX1 arr_reg_32__14_ ( .D(n4003), .CLK(clk), .Q(arr[526]) );
  DFFPOSX1 arr_reg_32__13_ ( .D(n4002), .CLK(clk), .Q(arr[525]) );
  DFFPOSX1 arr_reg_32__12_ ( .D(n4001), .CLK(clk), .Q(arr[524]) );
  DFFPOSX1 arr_reg_32__11_ ( .D(n4000), .CLK(clk), .Q(arr[523]) );
  DFFPOSX1 arr_reg_32__10_ ( .D(n3999), .CLK(clk), .Q(arr[522]) );
  DFFPOSX1 arr_reg_32__9_ ( .D(n3998), .CLK(clk), .Q(arr[521]) );
  DFFPOSX1 arr_reg_32__8_ ( .D(n3997), .CLK(clk), .Q(arr[520]) );
  DFFPOSX1 arr_reg_32__7_ ( .D(n3996), .CLK(clk), .Q(arr[519]) );
  DFFPOSX1 arr_reg_32__6_ ( .D(n3995), .CLK(clk), .Q(arr[518]) );
  DFFPOSX1 arr_reg_32__5_ ( .D(n3994), .CLK(clk), .Q(arr[517]) );
  DFFPOSX1 arr_reg_32__4_ ( .D(n3993), .CLK(clk), .Q(arr[516]) );
  DFFPOSX1 arr_reg_32__3_ ( .D(n3992), .CLK(clk), .Q(arr[515]) );
  DFFPOSX1 arr_reg_32__2_ ( .D(n3991), .CLK(clk), .Q(arr[514]) );
  DFFPOSX1 arr_reg_32__1_ ( .D(n3990), .CLK(clk), .Q(arr[513]) );
  DFFPOSX1 arr_reg_32__0_ ( .D(n3989), .CLK(clk), .Q(arr[512]) );
  DFFPOSX1 arr_reg_31__15_ ( .D(n3988), .CLK(clk), .Q(arr[511]) );
  DFFPOSX1 arr_reg_31__14_ ( .D(n3987), .CLK(clk), .Q(arr[510]) );
  DFFPOSX1 arr_reg_31__13_ ( .D(n3986), .CLK(clk), .Q(arr[509]) );
  DFFPOSX1 arr_reg_31__12_ ( .D(n3985), .CLK(clk), .Q(arr[508]) );
  DFFPOSX1 arr_reg_31__11_ ( .D(n3984), .CLK(clk), .Q(arr[507]) );
  DFFPOSX1 arr_reg_31__10_ ( .D(n3983), .CLK(clk), .Q(arr[506]) );
  DFFPOSX1 arr_reg_31__9_ ( .D(n3982), .CLK(clk), .Q(arr[505]) );
  DFFPOSX1 arr_reg_31__8_ ( .D(n3981), .CLK(clk), .Q(arr[504]) );
  DFFPOSX1 arr_reg_31__7_ ( .D(n3980), .CLK(clk), .Q(arr[503]) );
  DFFPOSX1 arr_reg_31__6_ ( .D(n3979), .CLK(clk), .Q(arr[502]) );
  DFFPOSX1 arr_reg_31__5_ ( .D(n3978), .CLK(clk), .Q(arr[501]) );
  DFFPOSX1 arr_reg_31__4_ ( .D(n3977), .CLK(clk), .Q(arr[500]) );
  DFFPOSX1 arr_reg_31__3_ ( .D(n3976), .CLK(clk), .Q(arr[499]) );
  DFFPOSX1 arr_reg_31__2_ ( .D(n3975), .CLK(clk), .Q(arr[498]) );
  DFFPOSX1 arr_reg_31__1_ ( .D(n3974), .CLK(clk), .Q(arr[497]) );
  DFFPOSX1 arr_reg_31__0_ ( .D(n3973), .CLK(clk), .Q(arr[496]) );
  DFFPOSX1 arr_reg_30__15_ ( .D(n3972), .CLK(clk), .Q(arr[495]) );
  DFFPOSX1 arr_reg_30__14_ ( .D(n3971), .CLK(clk), .Q(arr[494]) );
  DFFPOSX1 arr_reg_30__13_ ( .D(n3970), .CLK(clk), .Q(arr[493]) );
  DFFPOSX1 arr_reg_30__12_ ( .D(n3969), .CLK(clk), .Q(arr[492]) );
  DFFPOSX1 arr_reg_30__11_ ( .D(n3968), .CLK(clk), .Q(arr[491]) );
  DFFPOSX1 arr_reg_30__10_ ( .D(n3967), .CLK(clk), .Q(arr[490]) );
  DFFPOSX1 arr_reg_30__9_ ( .D(n3966), .CLK(clk), .Q(arr[489]) );
  DFFPOSX1 arr_reg_30__8_ ( .D(n3965), .CLK(clk), .Q(arr[488]) );
  DFFPOSX1 arr_reg_30__7_ ( .D(n3964), .CLK(clk), .Q(arr[487]) );
  DFFPOSX1 arr_reg_30__6_ ( .D(n3963), .CLK(clk), .Q(arr[486]) );
  DFFPOSX1 arr_reg_30__5_ ( .D(n3962), .CLK(clk), .Q(arr[485]) );
  DFFPOSX1 arr_reg_30__4_ ( .D(n3961), .CLK(clk), .Q(arr[484]) );
  DFFPOSX1 arr_reg_30__3_ ( .D(n3960), .CLK(clk), .Q(arr[483]) );
  DFFPOSX1 arr_reg_30__2_ ( .D(n3959), .CLK(clk), .Q(arr[482]) );
  DFFPOSX1 arr_reg_30__1_ ( .D(n3958), .CLK(clk), .Q(arr[481]) );
  DFFPOSX1 arr_reg_30__0_ ( .D(n3957), .CLK(clk), .Q(arr[480]) );
  DFFPOSX1 arr_reg_29__15_ ( .D(n3956), .CLK(clk), .Q(arr[479]) );
  DFFPOSX1 arr_reg_29__14_ ( .D(n3955), .CLK(clk), .Q(arr[478]) );
  DFFPOSX1 arr_reg_29__13_ ( .D(n3954), .CLK(clk), .Q(arr[477]) );
  DFFPOSX1 arr_reg_29__12_ ( .D(n3953), .CLK(clk), .Q(arr[476]) );
  DFFPOSX1 arr_reg_29__11_ ( .D(n3952), .CLK(clk), .Q(arr[475]) );
  DFFPOSX1 arr_reg_29__10_ ( .D(n3951), .CLK(clk), .Q(arr[474]) );
  DFFPOSX1 arr_reg_29__9_ ( .D(n3950), .CLK(clk), .Q(arr[473]) );
  DFFPOSX1 arr_reg_29__8_ ( .D(n3949), .CLK(clk), .Q(arr[472]) );
  DFFPOSX1 arr_reg_29__7_ ( .D(n3948), .CLK(clk), .Q(arr[471]) );
  DFFPOSX1 arr_reg_29__6_ ( .D(n3947), .CLK(clk), .Q(arr[470]) );
  DFFPOSX1 arr_reg_29__5_ ( .D(n3946), .CLK(clk), .Q(arr[469]) );
  DFFPOSX1 arr_reg_29__4_ ( .D(n3945), .CLK(clk), .Q(arr[468]) );
  DFFPOSX1 arr_reg_29__3_ ( .D(n3944), .CLK(clk), .Q(arr[467]) );
  DFFPOSX1 arr_reg_29__2_ ( .D(n3943), .CLK(clk), .Q(arr[466]) );
  DFFPOSX1 arr_reg_29__1_ ( .D(n3942), .CLK(clk), .Q(arr[465]) );
  DFFPOSX1 arr_reg_29__0_ ( .D(n3941), .CLK(clk), .Q(arr[464]) );
  DFFPOSX1 arr_reg_28__15_ ( .D(n3940), .CLK(clk), .Q(arr[463]) );
  DFFPOSX1 arr_reg_28__14_ ( .D(n3939), .CLK(clk), .Q(arr[462]) );
  DFFPOSX1 arr_reg_28__13_ ( .D(n3938), .CLK(clk), .Q(arr[461]) );
  DFFPOSX1 arr_reg_28__12_ ( .D(n3937), .CLK(clk), .Q(arr[460]) );
  DFFPOSX1 arr_reg_28__11_ ( .D(n3936), .CLK(clk), .Q(arr[459]) );
  DFFPOSX1 arr_reg_28__10_ ( .D(n3935), .CLK(clk), .Q(arr[458]) );
  DFFPOSX1 arr_reg_28__9_ ( .D(n3934), .CLK(clk), .Q(arr[457]) );
  DFFPOSX1 arr_reg_28__8_ ( .D(n3933), .CLK(clk), .Q(arr[456]) );
  DFFPOSX1 arr_reg_28__7_ ( .D(n3932), .CLK(clk), .Q(arr[455]) );
  DFFPOSX1 arr_reg_28__6_ ( .D(n3931), .CLK(clk), .Q(arr[454]) );
  DFFPOSX1 arr_reg_28__5_ ( .D(n3930), .CLK(clk), .Q(arr[453]) );
  DFFPOSX1 arr_reg_28__4_ ( .D(n3929), .CLK(clk), .Q(arr[452]) );
  DFFPOSX1 arr_reg_28__3_ ( .D(n3928), .CLK(clk), .Q(arr[451]) );
  DFFPOSX1 arr_reg_28__2_ ( .D(n3927), .CLK(clk), .Q(arr[450]) );
  DFFPOSX1 arr_reg_28__1_ ( .D(n3926), .CLK(clk), .Q(arr[449]) );
  DFFPOSX1 arr_reg_28__0_ ( .D(n3925), .CLK(clk), .Q(arr[448]) );
  DFFPOSX1 arr_reg_27__15_ ( .D(n3924), .CLK(clk), .Q(arr[447]) );
  DFFPOSX1 arr_reg_27__14_ ( .D(n3923), .CLK(clk), .Q(arr[446]) );
  DFFPOSX1 arr_reg_27__13_ ( .D(n3922), .CLK(clk), .Q(arr[445]) );
  DFFPOSX1 arr_reg_27__12_ ( .D(n3921), .CLK(clk), .Q(arr[444]) );
  DFFPOSX1 arr_reg_27__11_ ( .D(n3920), .CLK(clk), .Q(arr[443]) );
  DFFPOSX1 arr_reg_27__10_ ( .D(n3919), .CLK(clk), .Q(arr[442]) );
  DFFPOSX1 arr_reg_27__9_ ( .D(n3918), .CLK(clk), .Q(arr[441]) );
  DFFPOSX1 arr_reg_27__8_ ( .D(n3917), .CLK(clk), .Q(arr[440]) );
  DFFPOSX1 arr_reg_27__7_ ( .D(n3916), .CLK(clk), .Q(arr[439]) );
  DFFPOSX1 arr_reg_27__6_ ( .D(n3915), .CLK(clk), .Q(arr[438]) );
  DFFPOSX1 arr_reg_27__5_ ( .D(n3914), .CLK(clk), .Q(arr[437]) );
  DFFPOSX1 arr_reg_27__4_ ( .D(n3913), .CLK(clk), .Q(arr[436]) );
  DFFPOSX1 arr_reg_27__3_ ( .D(n3912), .CLK(clk), .Q(arr[435]) );
  DFFPOSX1 arr_reg_27__2_ ( .D(n3911), .CLK(clk), .Q(arr[434]) );
  DFFPOSX1 arr_reg_27__1_ ( .D(n3910), .CLK(clk), .Q(arr[433]) );
  DFFPOSX1 arr_reg_27__0_ ( .D(n3909), .CLK(clk), .Q(arr[432]) );
  DFFPOSX1 arr_reg_26__15_ ( .D(n3908), .CLK(clk), .Q(arr[431]) );
  DFFPOSX1 arr_reg_26__14_ ( .D(n3907), .CLK(clk), .Q(arr[430]) );
  DFFPOSX1 arr_reg_26__13_ ( .D(n3906), .CLK(clk), .Q(arr[429]) );
  DFFPOSX1 arr_reg_26__12_ ( .D(n3905), .CLK(clk), .Q(arr[428]) );
  DFFPOSX1 arr_reg_26__11_ ( .D(n3904), .CLK(clk), .Q(arr[427]) );
  DFFPOSX1 arr_reg_26__10_ ( .D(n3903), .CLK(clk), .Q(arr[426]) );
  DFFPOSX1 arr_reg_26__9_ ( .D(n3902), .CLK(clk), .Q(arr[425]) );
  DFFPOSX1 arr_reg_26__8_ ( .D(n3901), .CLK(clk), .Q(arr[424]) );
  DFFPOSX1 arr_reg_26__7_ ( .D(n3900), .CLK(clk), .Q(arr[423]) );
  DFFPOSX1 arr_reg_26__6_ ( .D(n3899), .CLK(clk), .Q(arr[422]) );
  DFFPOSX1 arr_reg_26__5_ ( .D(n3898), .CLK(clk), .Q(arr[421]) );
  DFFPOSX1 arr_reg_26__4_ ( .D(n3897), .CLK(clk), .Q(arr[420]) );
  DFFPOSX1 arr_reg_26__3_ ( .D(n3896), .CLK(clk), .Q(arr[419]) );
  DFFPOSX1 arr_reg_26__2_ ( .D(n3895), .CLK(clk), .Q(arr[418]) );
  DFFPOSX1 arr_reg_26__1_ ( .D(n3894), .CLK(clk), .Q(arr[417]) );
  DFFPOSX1 arr_reg_26__0_ ( .D(n3893), .CLK(clk), .Q(arr[416]) );
  DFFPOSX1 arr_reg_25__15_ ( .D(n3892), .CLK(clk), .Q(arr[415]) );
  DFFPOSX1 arr_reg_25__14_ ( .D(n3891), .CLK(clk), .Q(arr[414]) );
  DFFPOSX1 arr_reg_25__13_ ( .D(n3890), .CLK(clk), .Q(arr[413]) );
  DFFPOSX1 arr_reg_25__12_ ( .D(n3889), .CLK(clk), .Q(arr[412]) );
  DFFPOSX1 arr_reg_25__11_ ( .D(n3888), .CLK(clk), .Q(arr[411]) );
  DFFPOSX1 arr_reg_25__10_ ( .D(n3887), .CLK(clk), .Q(arr[410]) );
  DFFPOSX1 arr_reg_25__9_ ( .D(n3886), .CLK(clk), .Q(arr[409]) );
  DFFPOSX1 arr_reg_25__8_ ( .D(n3885), .CLK(clk), .Q(arr[408]) );
  DFFPOSX1 arr_reg_25__7_ ( .D(n3884), .CLK(clk), .Q(arr[407]) );
  DFFPOSX1 arr_reg_25__6_ ( .D(n3883), .CLK(clk), .Q(arr[406]) );
  DFFPOSX1 arr_reg_25__5_ ( .D(n3882), .CLK(clk), .Q(arr[405]) );
  DFFPOSX1 arr_reg_25__4_ ( .D(n3881), .CLK(clk), .Q(arr[404]) );
  DFFPOSX1 arr_reg_25__3_ ( .D(n3880), .CLK(clk), .Q(arr[403]) );
  DFFPOSX1 arr_reg_25__2_ ( .D(n3879), .CLK(clk), .Q(arr[402]) );
  DFFPOSX1 arr_reg_25__1_ ( .D(n3878), .CLK(clk), .Q(arr[401]) );
  DFFPOSX1 arr_reg_25__0_ ( .D(n3877), .CLK(clk), .Q(arr[400]) );
  DFFPOSX1 arr_reg_24__15_ ( .D(n3876), .CLK(clk), .Q(arr[399]) );
  DFFPOSX1 arr_reg_24__14_ ( .D(n3875), .CLK(clk), .Q(arr[398]) );
  DFFPOSX1 arr_reg_24__13_ ( .D(n3874), .CLK(clk), .Q(arr[397]) );
  DFFPOSX1 arr_reg_24__12_ ( .D(n3873), .CLK(clk), .Q(arr[396]) );
  DFFPOSX1 arr_reg_24__11_ ( .D(n3872), .CLK(clk), .Q(arr[395]) );
  DFFPOSX1 arr_reg_24__10_ ( .D(n3871), .CLK(clk), .Q(arr[394]) );
  DFFPOSX1 arr_reg_24__9_ ( .D(n3870), .CLK(clk), .Q(arr[393]) );
  DFFPOSX1 arr_reg_24__8_ ( .D(n3869), .CLK(clk), .Q(arr[392]) );
  DFFPOSX1 arr_reg_24__7_ ( .D(n3868), .CLK(clk), .Q(arr[391]) );
  DFFPOSX1 arr_reg_24__6_ ( .D(n3867), .CLK(clk), .Q(arr[390]) );
  DFFPOSX1 arr_reg_24__5_ ( .D(n3866), .CLK(clk), .Q(arr[389]) );
  DFFPOSX1 arr_reg_24__4_ ( .D(n3865), .CLK(clk), .Q(arr[388]) );
  DFFPOSX1 arr_reg_24__3_ ( .D(n3864), .CLK(clk), .Q(arr[387]) );
  DFFPOSX1 arr_reg_24__2_ ( .D(n3863), .CLK(clk), .Q(arr[386]) );
  DFFPOSX1 arr_reg_24__1_ ( .D(n3862), .CLK(clk), .Q(arr[385]) );
  DFFPOSX1 arr_reg_24__0_ ( .D(n3861), .CLK(clk), .Q(arr[384]) );
  DFFPOSX1 arr_reg_23__15_ ( .D(n3860), .CLK(clk), .Q(arr[383]) );
  DFFPOSX1 arr_reg_23__14_ ( .D(n3859), .CLK(clk), .Q(arr[382]) );
  DFFPOSX1 arr_reg_23__13_ ( .D(n3858), .CLK(clk), .Q(arr[381]) );
  DFFPOSX1 arr_reg_23__12_ ( .D(n3857), .CLK(clk), .Q(arr[380]) );
  DFFPOSX1 arr_reg_23__11_ ( .D(n3856), .CLK(clk), .Q(arr[379]) );
  DFFPOSX1 arr_reg_23__10_ ( .D(n3855), .CLK(clk), .Q(arr[378]) );
  DFFPOSX1 arr_reg_23__9_ ( .D(n3854), .CLK(clk), .Q(arr[377]) );
  DFFPOSX1 arr_reg_23__8_ ( .D(n3853), .CLK(clk), .Q(arr[376]) );
  DFFPOSX1 arr_reg_23__7_ ( .D(n3852), .CLK(clk), .Q(arr[375]) );
  DFFPOSX1 arr_reg_23__6_ ( .D(n3851), .CLK(clk), .Q(arr[374]) );
  DFFPOSX1 arr_reg_23__5_ ( .D(n3850), .CLK(clk), .Q(arr[373]) );
  DFFPOSX1 arr_reg_23__4_ ( .D(n3849), .CLK(clk), .Q(arr[372]) );
  DFFPOSX1 arr_reg_23__3_ ( .D(n3848), .CLK(clk), .Q(arr[371]) );
  DFFPOSX1 arr_reg_23__2_ ( .D(n3847), .CLK(clk), .Q(arr[370]) );
  DFFPOSX1 arr_reg_23__1_ ( .D(n3846), .CLK(clk), .Q(arr[369]) );
  DFFPOSX1 arr_reg_23__0_ ( .D(n3845), .CLK(clk), .Q(arr[368]) );
  DFFPOSX1 arr_reg_22__15_ ( .D(n3844), .CLK(clk), .Q(arr[367]) );
  DFFPOSX1 arr_reg_22__14_ ( .D(n3843), .CLK(clk), .Q(arr[366]) );
  DFFPOSX1 arr_reg_22__13_ ( .D(n3842), .CLK(clk), .Q(arr[365]) );
  DFFPOSX1 arr_reg_22__12_ ( .D(n3841), .CLK(clk), .Q(arr[364]) );
  DFFPOSX1 arr_reg_22__11_ ( .D(n3840), .CLK(clk), .Q(arr[363]) );
  DFFPOSX1 arr_reg_22__10_ ( .D(n3839), .CLK(clk), .Q(arr[362]) );
  DFFPOSX1 arr_reg_22__9_ ( .D(n3838), .CLK(clk), .Q(arr[361]) );
  DFFPOSX1 arr_reg_22__8_ ( .D(n3837), .CLK(clk), .Q(arr[360]) );
  DFFPOSX1 arr_reg_22__7_ ( .D(n3836), .CLK(clk), .Q(arr[359]) );
  DFFPOSX1 arr_reg_22__6_ ( .D(n3835), .CLK(clk), .Q(arr[358]) );
  DFFPOSX1 arr_reg_22__5_ ( .D(n3834), .CLK(clk), .Q(arr[357]) );
  DFFPOSX1 arr_reg_22__4_ ( .D(n3833), .CLK(clk), .Q(arr[356]) );
  DFFPOSX1 arr_reg_22__3_ ( .D(n3832), .CLK(clk), .Q(arr[355]) );
  DFFPOSX1 arr_reg_22__2_ ( .D(n3831), .CLK(clk), .Q(arr[354]) );
  DFFPOSX1 arr_reg_22__1_ ( .D(n3830), .CLK(clk), .Q(arr[353]) );
  DFFPOSX1 arr_reg_22__0_ ( .D(n3829), .CLK(clk), .Q(arr[352]) );
  DFFPOSX1 arr_reg_21__15_ ( .D(n3828), .CLK(clk), .Q(arr[351]) );
  DFFPOSX1 arr_reg_21__14_ ( .D(n3827), .CLK(clk), .Q(arr[350]) );
  DFFPOSX1 arr_reg_21__13_ ( .D(n3826), .CLK(clk), .Q(arr[349]) );
  DFFPOSX1 arr_reg_21__12_ ( .D(n3825), .CLK(clk), .Q(arr[348]) );
  DFFPOSX1 arr_reg_21__11_ ( .D(n3824), .CLK(clk), .Q(arr[347]) );
  DFFPOSX1 arr_reg_21__10_ ( .D(n3823), .CLK(clk), .Q(arr[346]) );
  DFFPOSX1 arr_reg_21__9_ ( .D(n3822), .CLK(clk), .Q(arr[345]) );
  DFFPOSX1 arr_reg_21__8_ ( .D(n3821), .CLK(clk), .Q(arr[344]) );
  DFFPOSX1 arr_reg_21__7_ ( .D(n3820), .CLK(clk), .Q(arr[343]) );
  DFFPOSX1 arr_reg_21__6_ ( .D(n3819), .CLK(clk), .Q(arr[342]) );
  DFFPOSX1 arr_reg_21__5_ ( .D(n3818), .CLK(clk), .Q(arr[341]) );
  DFFPOSX1 arr_reg_21__4_ ( .D(n3817), .CLK(clk), .Q(arr[340]) );
  DFFPOSX1 arr_reg_21__3_ ( .D(n3816), .CLK(clk), .Q(arr[339]) );
  DFFPOSX1 arr_reg_21__2_ ( .D(n3815), .CLK(clk), .Q(arr[338]) );
  DFFPOSX1 arr_reg_21__1_ ( .D(n3814), .CLK(clk), .Q(arr[337]) );
  DFFPOSX1 arr_reg_21__0_ ( .D(n3813), .CLK(clk), .Q(arr[336]) );
  DFFPOSX1 arr_reg_20__15_ ( .D(n3812), .CLK(clk), .Q(arr[335]) );
  DFFPOSX1 arr_reg_20__14_ ( .D(n3811), .CLK(clk), .Q(arr[334]) );
  DFFPOSX1 arr_reg_20__13_ ( .D(n3810), .CLK(clk), .Q(arr[333]) );
  DFFPOSX1 arr_reg_20__12_ ( .D(n3809), .CLK(clk), .Q(arr[332]) );
  DFFPOSX1 arr_reg_20__11_ ( .D(n3808), .CLK(clk), .Q(arr[331]) );
  DFFPOSX1 arr_reg_20__10_ ( .D(n3807), .CLK(clk), .Q(arr[330]) );
  DFFPOSX1 arr_reg_20__9_ ( .D(n3806), .CLK(clk), .Q(arr[329]) );
  DFFPOSX1 arr_reg_20__8_ ( .D(n3805), .CLK(clk), .Q(arr[328]) );
  DFFPOSX1 arr_reg_20__7_ ( .D(n3804), .CLK(clk), .Q(arr[327]) );
  DFFPOSX1 arr_reg_20__6_ ( .D(n3803), .CLK(clk), .Q(arr[326]) );
  DFFPOSX1 arr_reg_20__5_ ( .D(n3802), .CLK(clk), .Q(arr[325]) );
  DFFPOSX1 arr_reg_20__4_ ( .D(n3801), .CLK(clk), .Q(arr[324]) );
  DFFPOSX1 arr_reg_20__3_ ( .D(n3800), .CLK(clk), .Q(arr[323]) );
  DFFPOSX1 arr_reg_20__2_ ( .D(n3799), .CLK(clk), .Q(arr[322]) );
  DFFPOSX1 arr_reg_20__1_ ( .D(n3798), .CLK(clk), .Q(arr[321]) );
  DFFPOSX1 arr_reg_20__0_ ( .D(n3797), .CLK(clk), .Q(arr[320]) );
  DFFPOSX1 arr_reg_19__15_ ( .D(n3796), .CLK(clk), .Q(arr[319]) );
  DFFPOSX1 arr_reg_19__14_ ( .D(n3795), .CLK(clk), .Q(arr[318]) );
  DFFPOSX1 arr_reg_19__13_ ( .D(n3794), .CLK(clk), .Q(arr[317]) );
  DFFPOSX1 arr_reg_19__12_ ( .D(n3793), .CLK(clk), .Q(arr[316]) );
  DFFPOSX1 arr_reg_19__11_ ( .D(n3792), .CLK(clk), .Q(arr[315]) );
  DFFPOSX1 arr_reg_19__10_ ( .D(n3791), .CLK(clk), .Q(arr[314]) );
  DFFPOSX1 arr_reg_19__9_ ( .D(n3790), .CLK(clk), .Q(arr[313]) );
  DFFPOSX1 arr_reg_19__8_ ( .D(n3789), .CLK(clk), .Q(arr[312]) );
  DFFPOSX1 arr_reg_19__7_ ( .D(n3788), .CLK(clk), .Q(arr[311]) );
  DFFPOSX1 arr_reg_19__6_ ( .D(n3787), .CLK(clk), .Q(arr[310]) );
  DFFPOSX1 arr_reg_19__5_ ( .D(n3786), .CLK(clk), .Q(arr[309]) );
  DFFPOSX1 arr_reg_19__4_ ( .D(n3785), .CLK(clk), .Q(arr[308]) );
  DFFPOSX1 arr_reg_19__3_ ( .D(n3784), .CLK(clk), .Q(arr[307]) );
  DFFPOSX1 arr_reg_19__2_ ( .D(n3783), .CLK(clk), .Q(arr[306]) );
  DFFPOSX1 arr_reg_19__1_ ( .D(n3782), .CLK(clk), .Q(arr[305]) );
  DFFPOSX1 arr_reg_19__0_ ( .D(n3781), .CLK(clk), .Q(arr[304]) );
  DFFPOSX1 arr_reg_18__15_ ( .D(n3780), .CLK(clk), .Q(arr[303]) );
  DFFPOSX1 arr_reg_18__14_ ( .D(n3779), .CLK(clk), .Q(arr[302]) );
  DFFPOSX1 arr_reg_18__13_ ( .D(n3778), .CLK(clk), .Q(arr[301]) );
  DFFPOSX1 arr_reg_18__12_ ( .D(n3777), .CLK(clk), .Q(arr[300]) );
  DFFPOSX1 arr_reg_18__11_ ( .D(n3776), .CLK(clk), .Q(arr[299]) );
  DFFPOSX1 arr_reg_18__10_ ( .D(n3775), .CLK(clk), .Q(arr[298]) );
  DFFPOSX1 arr_reg_18__9_ ( .D(n3774), .CLK(clk), .Q(arr[297]) );
  DFFPOSX1 arr_reg_18__8_ ( .D(n3773), .CLK(clk), .Q(arr[296]) );
  DFFPOSX1 arr_reg_18__7_ ( .D(n3772), .CLK(clk), .Q(arr[295]) );
  DFFPOSX1 arr_reg_18__6_ ( .D(n3771), .CLK(clk), .Q(arr[294]) );
  DFFPOSX1 arr_reg_18__5_ ( .D(n3770), .CLK(clk), .Q(arr[293]) );
  DFFPOSX1 arr_reg_18__4_ ( .D(n3769), .CLK(clk), .Q(arr[292]) );
  DFFPOSX1 arr_reg_18__3_ ( .D(n3768), .CLK(clk), .Q(arr[291]) );
  DFFPOSX1 arr_reg_18__2_ ( .D(n3767), .CLK(clk), .Q(arr[290]) );
  DFFPOSX1 arr_reg_18__1_ ( .D(n3766), .CLK(clk), .Q(arr[289]) );
  DFFPOSX1 arr_reg_18__0_ ( .D(n3765), .CLK(clk), .Q(arr[288]) );
  DFFPOSX1 arr_reg_17__15_ ( .D(n3764), .CLK(clk), .Q(arr[287]) );
  DFFPOSX1 arr_reg_17__14_ ( .D(n3763), .CLK(clk), .Q(arr[286]) );
  DFFPOSX1 arr_reg_17__13_ ( .D(n3762), .CLK(clk), .Q(arr[285]) );
  DFFPOSX1 arr_reg_17__12_ ( .D(n3761), .CLK(clk), .Q(arr[284]) );
  DFFPOSX1 arr_reg_17__11_ ( .D(n3760), .CLK(clk), .Q(arr[283]) );
  DFFPOSX1 arr_reg_17__10_ ( .D(n3759), .CLK(clk), .Q(arr[282]) );
  DFFPOSX1 arr_reg_17__9_ ( .D(n3758), .CLK(clk), .Q(arr[281]) );
  DFFPOSX1 arr_reg_17__8_ ( .D(n3757), .CLK(clk), .Q(arr[280]) );
  DFFPOSX1 arr_reg_17__7_ ( .D(n3756), .CLK(clk), .Q(arr[279]) );
  DFFPOSX1 arr_reg_17__6_ ( .D(n3755), .CLK(clk), .Q(arr[278]) );
  DFFPOSX1 arr_reg_17__5_ ( .D(n3754), .CLK(clk), .Q(arr[277]) );
  DFFPOSX1 arr_reg_17__4_ ( .D(n3753), .CLK(clk), .Q(arr[276]) );
  DFFPOSX1 arr_reg_17__3_ ( .D(n3752), .CLK(clk), .Q(arr[275]) );
  DFFPOSX1 arr_reg_17__2_ ( .D(n3751), .CLK(clk), .Q(arr[274]) );
  DFFPOSX1 arr_reg_17__1_ ( .D(n3750), .CLK(clk), .Q(arr[273]) );
  DFFPOSX1 arr_reg_17__0_ ( .D(n3749), .CLK(clk), .Q(arr[272]) );
  DFFPOSX1 arr_reg_16__15_ ( .D(n3748), .CLK(clk), .Q(arr[271]) );
  DFFPOSX1 arr_reg_16__14_ ( .D(n3747), .CLK(clk), .Q(arr[270]) );
  DFFPOSX1 arr_reg_16__13_ ( .D(n3746), .CLK(clk), .Q(arr[269]) );
  DFFPOSX1 arr_reg_16__12_ ( .D(n3745), .CLK(clk), .Q(arr[268]) );
  DFFPOSX1 arr_reg_16__11_ ( .D(n3744), .CLK(clk), .Q(arr[267]) );
  DFFPOSX1 arr_reg_16__10_ ( .D(n3743), .CLK(clk), .Q(arr[266]) );
  DFFPOSX1 arr_reg_16__9_ ( .D(n3742), .CLK(clk), .Q(arr[265]) );
  DFFPOSX1 arr_reg_16__8_ ( .D(n3741), .CLK(clk), .Q(arr[264]) );
  DFFPOSX1 arr_reg_16__7_ ( .D(n3740), .CLK(clk), .Q(arr[263]) );
  DFFPOSX1 arr_reg_16__6_ ( .D(n3739), .CLK(clk), .Q(arr[262]) );
  DFFPOSX1 arr_reg_16__5_ ( .D(n3738), .CLK(clk), .Q(arr[261]) );
  DFFPOSX1 arr_reg_16__4_ ( .D(n3737), .CLK(clk), .Q(arr[260]) );
  DFFPOSX1 arr_reg_16__3_ ( .D(n3736), .CLK(clk), .Q(arr[259]) );
  DFFPOSX1 arr_reg_16__2_ ( .D(n3735), .CLK(clk), .Q(arr[258]) );
  DFFPOSX1 arr_reg_16__1_ ( .D(n3734), .CLK(clk), .Q(arr[257]) );
  DFFPOSX1 arr_reg_16__0_ ( .D(n3733), .CLK(clk), .Q(arr[256]) );
  DFFPOSX1 arr_reg_15__15_ ( .D(n3732), .CLK(clk), .Q(arr[255]) );
  DFFPOSX1 arr_reg_15__14_ ( .D(n3731), .CLK(clk), .Q(arr[254]) );
  DFFPOSX1 arr_reg_15__13_ ( .D(n3730), .CLK(clk), .Q(arr[253]) );
  DFFPOSX1 arr_reg_15__12_ ( .D(n3729), .CLK(clk), .Q(arr[252]) );
  DFFPOSX1 arr_reg_15__11_ ( .D(n3728), .CLK(clk), .Q(arr[251]) );
  DFFPOSX1 arr_reg_15__10_ ( .D(n3727), .CLK(clk), .Q(arr[250]) );
  DFFPOSX1 arr_reg_15__9_ ( .D(n3726), .CLK(clk), .Q(arr[249]) );
  DFFPOSX1 arr_reg_15__8_ ( .D(n3725), .CLK(clk), .Q(arr[248]) );
  DFFPOSX1 arr_reg_15__7_ ( .D(n3724), .CLK(clk), .Q(arr[247]) );
  DFFPOSX1 arr_reg_15__6_ ( .D(n3723), .CLK(clk), .Q(arr[246]) );
  DFFPOSX1 arr_reg_15__5_ ( .D(n3722), .CLK(clk), .Q(arr[245]) );
  DFFPOSX1 arr_reg_15__4_ ( .D(n3721), .CLK(clk), .Q(arr[244]) );
  DFFPOSX1 arr_reg_15__3_ ( .D(n3720), .CLK(clk), .Q(arr[243]) );
  DFFPOSX1 arr_reg_15__2_ ( .D(n3719), .CLK(clk), .Q(arr[242]) );
  DFFPOSX1 arr_reg_15__1_ ( .D(n3718), .CLK(clk), .Q(arr[241]) );
  DFFPOSX1 arr_reg_15__0_ ( .D(n3717), .CLK(clk), .Q(arr[240]) );
  DFFPOSX1 arr_reg_14__15_ ( .D(n3716), .CLK(clk), .Q(arr[239]) );
  DFFPOSX1 arr_reg_14__14_ ( .D(n3715), .CLK(clk), .Q(arr[238]) );
  DFFPOSX1 arr_reg_14__13_ ( .D(n3714), .CLK(clk), .Q(arr[237]) );
  DFFPOSX1 arr_reg_14__12_ ( .D(n3713), .CLK(clk), .Q(arr[236]) );
  DFFPOSX1 arr_reg_14__11_ ( .D(n3712), .CLK(clk), .Q(arr[235]) );
  DFFPOSX1 arr_reg_14__10_ ( .D(n3711), .CLK(clk), .Q(arr[234]) );
  DFFPOSX1 arr_reg_14__9_ ( .D(n3710), .CLK(clk), .Q(arr[233]) );
  DFFPOSX1 arr_reg_14__8_ ( .D(n3709), .CLK(clk), .Q(arr[232]) );
  DFFPOSX1 arr_reg_14__7_ ( .D(n3708), .CLK(clk), .Q(arr[231]) );
  DFFPOSX1 arr_reg_14__6_ ( .D(n3707), .CLK(clk), .Q(arr[230]) );
  DFFPOSX1 arr_reg_14__5_ ( .D(n3706), .CLK(clk), .Q(arr[229]) );
  DFFPOSX1 arr_reg_14__4_ ( .D(n3705), .CLK(clk), .Q(arr[228]) );
  DFFPOSX1 arr_reg_14__3_ ( .D(n3704), .CLK(clk), .Q(arr[227]) );
  DFFPOSX1 arr_reg_14__2_ ( .D(n3703), .CLK(clk), .Q(arr[226]) );
  DFFPOSX1 arr_reg_14__1_ ( .D(n3702), .CLK(clk), .Q(arr[225]) );
  DFFPOSX1 arr_reg_14__0_ ( .D(n3701), .CLK(clk), .Q(arr[224]) );
  DFFPOSX1 arr_reg_13__15_ ( .D(n3700), .CLK(clk), .Q(arr[223]) );
  DFFPOSX1 arr_reg_13__14_ ( .D(n3699), .CLK(clk), .Q(arr[222]) );
  DFFPOSX1 arr_reg_13__13_ ( .D(n3698), .CLK(clk), .Q(arr[221]) );
  DFFPOSX1 arr_reg_13__12_ ( .D(n3697), .CLK(clk), .Q(arr[220]) );
  DFFPOSX1 arr_reg_13__11_ ( .D(n3696), .CLK(clk), .Q(arr[219]) );
  DFFPOSX1 arr_reg_13__10_ ( .D(n3695), .CLK(clk), .Q(arr[218]) );
  DFFPOSX1 arr_reg_13__9_ ( .D(n3694), .CLK(clk), .Q(arr[217]) );
  DFFPOSX1 arr_reg_13__8_ ( .D(n3693), .CLK(clk), .Q(arr[216]) );
  DFFPOSX1 arr_reg_13__7_ ( .D(n3692), .CLK(clk), .Q(arr[215]) );
  DFFPOSX1 arr_reg_13__6_ ( .D(n3691), .CLK(clk), .Q(arr[214]) );
  DFFPOSX1 arr_reg_13__5_ ( .D(n3690), .CLK(clk), .Q(arr[213]) );
  DFFPOSX1 arr_reg_13__4_ ( .D(n3689), .CLK(clk), .Q(arr[212]) );
  DFFPOSX1 arr_reg_13__3_ ( .D(n3688), .CLK(clk), .Q(arr[211]) );
  DFFPOSX1 arr_reg_13__2_ ( .D(n3687), .CLK(clk), .Q(arr[210]) );
  DFFPOSX1 arr_reg_13__1_ ( .D(n3686), .CLK(clk), .Q(arr[209]) );
  DFFPOSX1 arr_reg_13__0_ ( .D(n3685), .CLK(clk), .Q(arr[208]) );
  DFFPOSX1 arr_reg_12__15_ ( .D(n3684), .CLK(clk), .Q(arr[207]) );
  DFFPOSX1 arr_reg_12__14_ ( .D(n3683), .CLK(clk), .Q(arr[206]) );
  DFFPOSX1 arr_reg_12__13_ ( .D(n3682), .CLK(clk), .Q(arr[205]) );
  DFFPOSX1 arr_reg_12__12_ ( .D(n3681), .CLK(clk), .Q(arr[204]) );
  DFFPOSX1 arr_reg_12__11_ ( .D(n3680), .CLK(clk), .Q(arr[203]) );
  DFFPOSX1 arr_reg_12__10_ ( .D(n3679), .CLK(clk), .Q(arr[202]) );
  DFFPOSX1 arr_reg_12__9_ ( .D(n3678), .CLK(clk), .Q(arr[201]) );
  DFFPOSX1 arr_reg_12__8_ ( .D(n3677), .CLK(clk), .Q(arr[200]) );
  DFFPOSX1 arr_reg_12__7_ ( .D(n3676), .CLK(clk), .Q(arr[199]) );
  DFFPOSX1 arr_reg_12__6_ ( .D(n3675), .CLK(clk), .Q(arr[198]) );
  DFFPOSX1 arr_reg_12__5_ ( .D(n3674), .CLK(clk), .Q(arr[197]) );
  DFFPOSX1 arr_reg_12__4_ ( .D(n3673), .CLK(clk), .Q(arr[196]) );
  DFFPOSX1 arr_reg_12__3_ ( .D(n3672), .CLK(clk), .Q(arr[195]) );
  DFFPOSX1 arr_reg_12__2_ ( .D(n3671), .CLK(clk), .Q(arr[194]) );
  DFFPOSX1 arr_reg_12__1_ ( .D(n3670), .CLK(clk), .Q(arr[193]) );
  DFFPOSX1 arr_reg_12__0_ ( .D(n3669), .CLK(clk), .Q(arr[192]) );
  DFFPOSX1 arr_reg_11__15_ ( .D(n3668), .CLK(clk), .Q(arr[191]) );
  DFFPOSX1 arr_reg_11__14_ ( .D(n3667), .CLK(clk), .Q(arr[190]) );
  DFFPOSX1 arr_reg_11__13_ ( .D(n3666), .CLK(clk), .Q(arr[189]) );
  DFFPOSX1 arr_reg_11__12_ ( .D(n3665), .CLK(clk), .Q(arr[188]) );
  DFFPOSX1 arr_reg_11__11_ ( .D(n3664), .CLK(clk), .Q(arr[187]) );
  DFFPOSX1 arr_reg_11__10_ ( .D(n3663), .CLK(clk), .Q(arr[186]) );
  DFFPOSX1 arr_reg_11__9_ ( .D(n3662), .CLK(clk), .Q(arr[185]) );
  DFFPOSX1 arr_reg_11__8_ ( .D(n3661), .CLK(clk), .Q(arr[184]) );
  DFFPOSX1 arr_reg_11__7_ ( .D(n3660), .CLK(clk), .Q(arr[183]) );
  DFFPOSX1 arr_reg_11__6_ ( .D(n3659), .CLK(clk), .Q(arr[182]) );
  DFFPOSX1 arr_reg_11__5_ ( .D(n3658), .CLK(clk), .Q(arr[181]) );
  DFFPOSX1 arr_reg_11__4_ ( .D(n3657), .CLK(clk), .Q(arr[180]) );
  DFFPOSX1 arr_reg_11__3_ ( .D(n3656), .CLK(clk), .Q(arr[179]) );
  DFFPOSX1 arr_reg_11__2_ ( .D(n3655), .CLK(clk), .Q(arr[178]) );
  DFFPOSX1 arr_reg_11__1_ ( .D(n3654), .CLK(clk), .Q(arr[177]) );
  DFFPOSX1 arr_reg_11__0_ ( .D(n3653), .CLK(clk), .Q(arr[176]) );
  DFFPOSX1 arr_reg_10__15_ ( .D(n3652), .CLK(clk), .Q(arr[175]) );
  DFFPOSX1 arr_reg_10__14_ ( .D(n3651), .CLK(clk), .Q(arr[174]) );
  DFFPOSX1 arr_reg_10__13_ ( .D(n3650), .CLK(clk), .Q(arr[173]) );
  DFFPOSX1 arr_reg_10__12_ ( .D(n3649), .CLK(clk), .Q(arr[172]) );
  DFFPOSX1 arr_reg_10__11_ ( .D(n3648), .CLK(clk), .Q(arr[171]) );
  DFFPOSX1 arr_reg_10__10_ ( .D(n3647), .CLK(clk), .Q(arr[170]) );
  DFFPOSX1 arr_reg_10__9_ ( .D(n3646), .CLK(clk), .Q(arr[169]) );
  DFFPOSX1 arr_reg_10__8_ ( .D(n3645), .CLK(clk), .Q(arr[168]) );
  DFFPOSX1 arr_reg_10__7_ ( .D(n3644), .CLK(clk), .Q(arr[167]) );
  DFFPOSX1 arr_reg_10__6_ ( .D(n3643), .CLK(clk), .Q(arr[166]) );
  DFFPOSX1 arr_reg_10__5_ ( .D(n3642), .CLK(clk), .Q(arr[165]) );
  DFFPOSX1 arr_reg_10__4_ ( .D(n3641), .CLK(clk), .Q(arr[164]) );
  DFFPOSX1 arr_reg_10__3_ ( .D(n3640), .CLK(clk), .Q(arr[163]) );
  DFFPOSX1 arr_reg_10__2_ ( .D(n3639), .CLK(clk), .Q(arr[162]) );
  DFFPOSX1 arr_reg_10__1_ ( .D(n3638), .CLK(clk), .Q(arr[161]) );
  DFFPOSX1 arr_reg_10__0_ ( .D(n3637), .CLK(clk), .Q(arr[160]) );
  DFFPOSX1 arr_reg_9__15_ ( .D(n3636), .CLK(clk), .Q(arr[159]) );
  DFFPOSX1 arr_reg_9__14_ ( .D(n3635), .CLK(clk), .Q(arr[158]) );
  DFFPOSX1 arr_reg_9__13_ ( .D(n3634), .CLK(clk), .Q(arr[157]) );
  DFFPOSX1 arr_reg_9__12_ ( .D(n3633), .CLK(clk), .Q(arr[156]) );
  DFFPOSX1 arr_reg_9__11_ ( .D(n3632), .CLK(clk), .Q(arr[155]) );
  DFFPOSX1 arr_reg_9__10_ ( .D(n3631), .CLK(clk), .Q(arr[154]) );
  DFFPOSX1 arr_reg_9__9_ ( .D(n3630), .CLK(clk), .Q(arr[153]) );
  DFFPOSX1 arr_reg_9__8_ ( .D(n3629), .CLK(clk), .Q(arr[152]) );
  DFFPOSX1 arr_reg_9__7_ ( .D(n3628), .CLK(clk), .Q(arr[151]) );
  DFFPOSX1 arr_reg_9__6_ ( .D(n3627), .CLK(clk), .Q(arr[150]) );
  DFFPOSX1 arr_reg_9__5_ ( .D(n3626), .CLK(clk), .Q(arr[149]) );
  DFFPOSX1 arr_reg_9__4_ ( .D(n3625), .CLK(clk), .Q(arr[148]) );
  DFFPOSX1 arr_reg_9__3_ ( .D(n3624), .CLK(clk), .Q(arr[147]) );
  DFFPOSX1 arr_reg_9__2_ ( .D(n3623), .CLK(clk), .Q(arr[146]) );
  DFFPOSX1 arr_reg_9__1_ ( .D(n3622), .CLK(clk), .Q(arr[145]) );
  DFFPOSX1 arr_reg_9__0_ ( .D(n3621), .CLK(clk), .Q(arr[144]) );
  DFFPOSX1 arr_reg_8__15_ ( .D(n3620), .CLK(clk), .Q(arr[143]) );
  DFFPOSX1 arr_reg_8__14_ ( .D(n3619), .CLK(clk), .Q(arr[142]) );
  DFFPOSX1 arr_reg_8__13_ ( .D(n3618), .CLK(clk), .Q(arr[141]) );
  DFFPOSX1 arr_reg_8__12_ ( .D(n3617), .CLK(clk), .Q(arr[140]) );
  DFFPOSX1 arr_reg_8__11_ ( .D(n3616), .CLK(clk), .Q(arr[139]) );
  DFFPOSX1 arr_reg_8__10_ ( .D(n3615), .CLK(clk), .Q(arr[138]) );
  DFFPOSX1 arr_reg_8__9_ ( .D(n3614), .CLK(clk), .Q(arr[137]) );
  DFFPOSX1 arr_reg_8__8_ ( .D(n3613), .CLK(clk), .Q(arr[136]) );
  DFFPOSX1 arr_reg_8__7_ ( .D(n3612), .CLK(clk), .Q(arr[135]) );
  DFFPOSX1 arr_reg_8__6_ ( .D(n3611), .CLK(clk), .Q(arr[134]) );
  DFFPOSX1 arr_reg_8__5_ ( .D(n3610), .CLK(clk), .Q(arr[133]) );
  DFFPOSX1 arr_reg_8__4_ ( .D(n3609), .CLK(clk), .Q(arr[132]) );
  DFFPOSX1 arr_reg_8__3_ ( .D(n3608), .CLK(clk), .Q(arr[131]) );
  DFFPOSX1 arr_reg_8__2_ ( .D(n3607), .CLK(clk), .Q(arr[130]) );
  DFFPOSX1 arr_reg_8__1_ ( .D(n3606), .CLK(clk), .Q(arr[129]) );
  DFFPOSX1 arr_reg_8__0_ ( .D(n3605), .CLK(clk), .Q(arr[128]) );
  DFFPOSX1 arr_reg_7__15_ ( .D(n3604), .CLK(clk), .Q(arr[127]) );
  DFFPOSX1 arr_reg_7__14_ ( .D(n3603), .CLK(clk), .Q(arr[126]) );
  DFFPOSX1 arr_reg_7__13_ ( .D(n3602), .CLK(clk), .Q(arr[125]) );
  DFFPOSX1 arr_reg_7__12_ ( .D(n3601), .CLK(clk), .Q(arr[124]) );
  DFFPOSX1 arr_reg_7__11_ ( .D(n3600), .CLK(clk), .Q(arr[123]) );
  DFFPOSX1 arr_reg_7__10_ ( .D(n3599), .CLK(clk), .Q(arr[122]) );
  DFFPOSX1 arr_reg_7__9_ ( .D(n3598), .CLK(clk), .Q(arr[121]) );
  DFFPOSX1 arr_reg_7__8_ ( .D(n3597), .CLK(clk), .Q(arr[120]) );
  DFFPOSX1 arr_reg_7__7_ ( .D(n3596), .CLK(clk), .Q(arr[119]) );
  DFFPOSX1 arr_reg_7__6_ ( .D(n3595), .CLK(clk), .Q(arr[118]) );
  DFFPOSX1 arr_reg_7__5_ ( .D(n3594), .CLK(clk), .Q(arr[117]) );
  DFFPOSX1 arr_reg_7__4_ ( .D(n3593), .CLK(clk), .Q(arr[116]) );
  DFFPOSX1 arr_reg_7__3_ ( .D(n3592), .CLK(clk), .Q(arr[115]) );
  DFFPOSX1 arr_reg_7__2_ ( .D(n3591), .CLK(clk), .Q(arr[114]) );
  DFFPOSX1 arr_reg_7__1_ ( .D(n3590), .CLK(clk), .Q(arr[113]) );
  DFFPOSX1 arr_reg_7__0_ ( .D(n3589), .CLK(clk), .Q(arr[112]) );
  DFFPOSX1 arr_reg_6__15_ ( .D(n3588), .CLK(clk), .Q(arr[111]) );
  DFFPOSX1 arr_reg_6__14_ ( .D(n3587), .CLK(clk), .Q(arr[110]) );
  DFFPOSX1 arr_reg_6__13_ ( .D(n3586), .CLK(clk), .Q(arr[109]) );
  DFFPOSX1 arr_reg_6__12_ ( .D(n3585), .CLK(clk), .Q(arr[108]) );
  DFFPOSX1 arr_reg_6__11_ ( .D(n3584), .CLK(clk), .Q(arr[107]) );
  DFFPOSX1 arr_reg_6__10_ ( .D(n3583), .CLK(clk), .Q(arr[106]) );
  DFFPOSX1 arr_reg_6__9_ ( .D(n3582), .CLK(clk), .Q(arr[105]) );
  DFFPOSX1 arr_reg_6__8_ ( .D(n3581), .CLK(clk), .Q(arr[104]) );
  DFFPOSX1 arr_reg_6__7_ ( .D(n3580), .CLK(clk), .Q(arr[103]) );
  DFFPOSX1 arr_reg_6__6_ ( .D(n3579), .CLK(clk), .Q(arr[102]) );
  DFFPOSX1 arr_reg_6__5_ ( .D(n3578), .CLK(clk), .Q(arr[101]) );
  DFFPOSX1 arr_reg_6__4_ ( .D(n3577), .CLK(clk), .Q(arr[100]) );
  DFFPOSX1 arr_reg_6__3_ ( .D(n3576), .CLK(clk), .Q(arr[99]) );
  DFFPOSX1 arr_reg_6__2_ ( .D(n3575), .CLK(clk), .Q(arr[98]) );
  DFFPOSX1 arr_reg_6__1_ ( .D(n3574), .CLK(clk), .Q(arr[97]) );
  DFFPOSX1 arr_reg_6__0_ ( .D(n3573), .CLK(clk), .Q(arr[96]) );
  DFFPOSX1 arr_reg_5__15_ ( .D(n3572), .CLK(clk), .Q(arr[95]) );
  DFFPOSX1 arr_reg_5__14_ ( .D(n3571), .CLK(clk), .Q(arr[94]) );
  DFFPOSX1 arr_reg_5__13_ ( .D(n3570), .CLK(clk), .Q(arr[93]) );
  DFFPOSX1 arr_reg_5__12_ ( .D(n3569), .CLK(clk), .Q(arr[92]) );
  DFFPOSX1 arr_reg_5__11_ ( .D(n3568), .CLK(clk), .Q(arr[91]) );
  DFFPOSX1 arr_reg_5__10_ ( .D(n3567), .CLK(clk), .Q(arr[90]) );
  DFFPOSX1 arr_reg_5__9_ ( .D(n3566), .CLK(clk), .Q(arr[89]) );
  DFFPOSX1 arr_reg_5__8_ ( .D(n3565), .CLK(clk), .Q(arr[88]) );
  DFFPOSX1 arr_reg_5__7_ ( .D(n3564), .CLK(clk), .Q(arr[87]) );
  DFFPOSX1 arr_reg_5__6_ ( .D(n3563), .CLK(clk), .Q(arr[86]) );
  DFFPOSX1 arr_reg_5__5_ ( .D(n3562), .CLK(clk), .Q(arr[85]) );
  DFFPOSX1 arr_reg_5__4_ ( .D(n3561), .CLK(clk), .Q(arr[84]) );
  DFFPOSX1 arr_reg_5__3_ ( .D(n3560), .CLK(clk), .Q(arr[83]) );
  DFFPOSX1 arr_reg_5__2_ ( .D(n3559), .CLK(clk), .Q(arr[82]) );
  DFFPOSX1 arr_reg_5__1_ ( .D(n3558), .CLK(clk), .Q(arr[81]) );
  DFFPOSX1 arr_reg_5__0_ ( .D(n3557), .CLK(clk), .Q(arr[80]) );
  DFFPOSX1 arr_reg_4__15_ ( .D(n3556), .CLK(clk), .Q(arr[79]) );
  DFFPOSX1 arr_reg_4__14_ ( .D(n3555), .CLK(clk), .Q(arr[78]) );
  DFFPOSX1 arr_reg_4__13_ ( .D(n3554), .CLK(clk), .Q(arr[77]) );
  DFFPOSX1 arr_reg_4__12_ ( .D(n3553), .CLK(clk), .Q(arr[76]) );
  DFFPOSX1 arr_reg_4__11_ ( .D(n3552), .CLK(clk), .Q(arr[75]) );
  DFFPOSX1 arr_reg_4__10_ ( .D(n3551), .CLK(clk), .Q(arr[74]) );
  DFFPOSX1 arr_reg_4__9_ ( .D(n3550), .CLK(clk), .Q(arr[73]) );
  DFFPOSX1 arr_reg_4__8_ ( .D(n3549), .CLK(clk), .Q(arr[72]) );
  DFFPOSX1 arr_reg_4__7_ ( .D(n3548), .CLK(clk), .Q(arr[71]) );
  DFFPOSX1 arr_reg_4__6_ ( .D(n3547), .CLK(clk), .Q(arr[70]) );
  DFFPOSX1 arr_reg_4__5_ ( .D(n3546), .CLK(clk), .Q(arr[69]) );
  DFFPOSX1 arr_reg_4__4_ ( .D(n3545), .CLK(clk), .Q(arr[68]) );
  DFFPOSX1 arr_reg_4__3_ ( .D(n3544), .CLK(clk), .Q(arr[67]) );
  DFFPOSX1 arr_reg_4__2_ ( .D(n3543), .CLK(clk), .Q(arr[66]) );
  DFFPOSX1 arr_reg_4__1_ ( .D(n3542), .CLK(clk), .Q(arr[65]) );
  DFFPOSX1 arr_reg_4__0_ ( .D(n3541), .CLK(clk), .Q(arr[64]) );
  DFFPOSX1 arr_reg_3__15_ ( .D(n3540), .CLK(clk), .Q(arr[63]) );
  DFFPOSX1 arr_reg_3__14_ ( .D(n3539), .CLK(clk), .Q(arr[62]) );
  DFFPOSX1 arr_reg_3__13_ ( .D(n3538), .CLK(clk), .Q(arr[61]) );
  DFFPOSX1 arr_reg_3__12_ ( .D(n3537), .CLK(clk), .Q(arr[60]) );
  DFFPOSX1 arr_reg_3__11_ ( .D(n3536), .CLK(clk), .Q(arr[59]) );
  DFFPOSX1 arr_reg_3__10_ ( .D(n3535), .CLK(clk), .Q(arr[58]) );
  DFFPOSX1 arr_reg_3__9_ ( .D(n3534), .CLK(clk), .Q(arr[57]) );
  DFFPOSX1 arr_reg_3__8_ ( .D(n3533), .CLK(clk), .Q(arr[56]) );
  DFFPOSX1 arr_reg_3__7_ ( .D(n3532), .CLK(clk), .Q(arr[55]) );
  DFFPOSX1 arr_reg_3__6_ ( .D(n3531), .CLK(clk), .Q(arr[54]) );
  DFFPOSX1 arr_reg_3__5_ ( .D(n3530), .CLK(clk), .Q(arr[53]) );
  DFFPOSX1 arr_reg_3__4_ ( .D(n3529), .CLK(clk), .Q(arr[52]) );
  DFFPOSX1 arr_reg_3__3_ ( .D(n3528), .CLK(clk), .Q(arr[51]) );
  DFFPOSX1 arr_reg_3__2_ ( .D(n3527), .CLK(clk), .Q(arr[50]) );
  DFFPOSX1 arr_reg_3__1_ ( .D(n3526), .CLK(clk), .Q(arr[49]) );
  DFFPOSX1 arr_reg_3__0_ ( .D(n3525), .CLK(clk), .Q(arr[48]) );
  DFFPOSX1 arr_reg_2__15_ ( .D(n3524), .CLK(clk), .Q(arr[47]) );
  DFFPOSX1 arr_reg_2__14_ ( .D(n3523), .CLK(clk), .Q(arr[46]) );
  DFFPOSX1 arr_reg_2__13_ ( .D(n3522), .CLK(clk), .Q(arr[45]) );
  DFFPOSX1 arr_reg_2__12_ ( .D(n3521), .CLK(clk), .Q(arr[44]) );
  DFFPOSX1 arr_reg_2__11_ ( .D(n3520), .CLK(clk), .Q(arr[43]) );
  DFFPOSX1 arr_reg_2__10_ ( .D(n3519), .CLK(clk), .Q(arr[42]) );
  DFFPOSX1 arr_reg_2__9_ ( .D(n3518), .CLK(clk), .Q(arr[41]) );
  DFFPOSX1 arr_reg_2__8_ ( .D(n3517), .CLK(clk), .Q(arr[40]) );
  DFFPOSX1 arr_reg_2__7_ ( .D(n3516), .CLK(clk), .Q(arr[39]) );
  DFFPOSX1 arr_reg_2__6_ ( .D(n3515), .CLK(clk), .Q(arr[38]) );
  DFFPOSX1 arr_reg_2__5_ ( .D(n3514), .CLK(clk), .Q(arr[37]) );
  DFFPOSX1 arr_reg_2__4_ ( .D(n3513), .CLK(clk), .Q(arr[36]) );
  DFFPOSX1 arr_reg_2__3_ ( .D(n3512), .CLK(clk), .Q(arr[35]) );
  DFFPOSX1 arr_reg_2__2_ ( .D(n3511), .CLK(clk), .Q(arr[34]) );
  DFFPOSX1 arr_reg_2__1_ ( .D(n3510), .CLK(clk), .Q(arr[33]) );
  DFFPOSX1 arr_reg_2__0_ ( .D(n3509), .CLK(clk), .Q(arr[32]) );
  DFFPOSX1 arr_reg_1__15_ ( .D(n3508), .CLK(clk), .Q(arr[31]) );
  DFFPOSX1 arr_reg_1__14_ ( .D(n3507), .CLK(clk), .Q(arr[30]) );
  DFFPOSX1 arr_reg_1__13_ ( .D(n3506), .CLK(clk), .Q(arr[29]) );
  DFFPOSX1 arr_reg_1__12_ ( .D(n3505), .CLK(clk), .Q(arr[28]) );
  DFFPOSX1 arr_reg_1__11_ ( .D(n3504), .CLK(clk), .Q(arr[27]) );
  DFFPOSX1 arr_reg_1__10_ ( .D(n3503), .CLK(clk), .Q(arr[26]) );
  DFFPOSX1 arr_reg_1__9_ ( .D(n3502), .CLK(clk), .Q(arr[25]) );
  DFFPOSX1 arr_reg_1__8_ ( .D(n3501), .CLK(clk), .Q(arr[24]) );
  DFFPOSX1 arr_reg_1__7_ ( .D(n3500), .CLK(clk), .Q(arr[23]) );
  DFFPOSX1 arr_reg_1__6_ ( .D(n3499), .CLK(clk), .Q(arr[22]) );
  DFFPOSX1 arr_reg_1__5_ ( .D(n3498), .CLK(clk), .Q(arr[21]) );
  DFFPOSX1 arr_reg_1__4_ ( .D(n3497), .CLK(clk), .Q(arr[20]) );
  DFFPOSX1 arr_reg_1__3_ ( .D(n3496), .CLK(clk), .Q(arr[19]) );
  DFFPOSX1 arr_reg_1__2_ ( .D(n3495), .CLK(clk), .Q(arr[18]) );
  DFFPOSX1 arr_reg_1__1_ ( .D(n3494), .CLK(clk), .Q(arr[17]) );
  DFFPOSX1 arr_reg_1__0_ ( .D(n3493), .CLK(clk), .Q(arr[16]) );
  DFFPOSX1 arr_reg_0__15_ ( .D(n3492), .CLK(clk), .Q(arr[15]) );
  DFFPOSX1 arr_reg_0__14_ ( .D(n3491), .CLK(clk), .Q(arr[14]) );
  DFFPOSX1 arr_reg_0__13_ ( .D(n3490), .CLK(clk), .Q(arr[13]) );
  DFFPOSX1 arr_reg_0__12_ ( .D(n3489), .CLK(clk), .Q(arr[12]) );
  DFFPOSX1 arr_reg_0__11_ ( .D(n3488), .CLK(clk), .Q(arr[11]) );
  DFFPOSX1 arr_reg_0__10_ ( .D(n3487), .CLK(clk), .Q(arr[10]) );
  DFFPOSX1 arr_reg_0__9_ ( .D(n3486), .CLK(clk), .Q(arr[9]) );
  DFFPOSX1 arr_reg_0__8_ ( .D(n3485), .CLK(clk), .Q(arr[8]) );
  DFFPOSX1 arr_reg_0__7_ ( .D(n3484), .CLK(clk), .Q(arr[7]) );
  DFFPOSX1 arr_reg_0__6_ ( .D(n3483), .CLK(clk), .Q(arr[6]) );
  DFFPOSX1 arr_reg_0__5_ ( .D(n3482), .CLK(clk), .Q(arr[5]) );
  DFFPOSX1 arr_reg_0__4_ ( .D(n3481), .CLK(clk), .Q(arr[4]) );
  DFFPOSX1 arr_reg_0__3_ ( .D(n3480), .CLK(clk), .Q(arr[3]) );
  DFFPOSX1 arr_reg_0__2_ ( .D(n3479), .CLK(clk), .Q(arr[2]) );
  DFFPOSX1 arr_reg_0__1_ ( .D(n3478), .CLK(clk), .Q(arr[1]) );
  DFFPOSX1 arr_reg_0__0_ ( .D(n3477), .CLK(clk), .Q(arr[0]) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n3476), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n3475), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n3474), .CLK(clk), .Q(n15) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n3473), .CLK(clk), .Q(n16) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n3472), .CLK(clk), .Q(n17) );
  DFFPOSX1 rd_ptr_reg_5_ ( .D(n3471), .CLK(clk), .Q(n18) );
  AOI22X1 U4 ( .A(n1130), .B(n2282), .C(n18), .D(n2283), .Y(n2281) );
  AOI22X1 U6 ( .A(n1129), .B(n2282), .C(n17), .D(n2283), .Y(n2284) );
  AOI22X1 U8 ( .A(n1128), .B(n2282), .C(n16), .D(n2283), .Y(n2285) );
  AOI22X1 U10 ( .A(n1127), .B(n2282), .C(n15), .D(n2283), .Y(n2286) );
  AOI22X1 U12 ( .A(n1126), .B(n2282), .C(n14), .D(n2283), .Y(n2287) );
  AOI22X1 U14 ( .A(n1125), .B(n2282), .C(n13), .D(n2283), .Y(n2288) );
  NOR2X1 U15 ( .A(n2283), .B(reset), .Y(n2282) );
  OAI21X1 U17 ( .A(n1336), .B(n1335), .C(n2292), .Y(n3477) );
  NAND2X1 U18 ( .A(arr[0]), .B(n1337), .Y(n2292) );
  OAI21X1 U19 ( .A(n1336), .B(n1334), .C(n2294), .Y(n3478) );
  NAND2X1 U20 ( .A(arr[1]), .B(n1336), .Y(n2294) );
  OAI21X1 U21 ( .A(n1336), .B(n1333), .C(n2296), .Y(n3479) );
  NAND2X1 U22 ( .A(arr[2]), .B(n1336), .Y(n2296) );
  OAI21X1 U23 ( .A(n1336), .B(n1332), .C(n2298), .Y(n3480) );
  NAND2X1 U24 ( .A(arr[3]), .B(n1337), .Y(n2298) );
  OAI21X1 U25 ( .A(n1336), .B(n1331), .C(n2300), .Y(n3481) );
  NAND2X1 U26 ( .A(arr[4]), .B(n1337), .Y(n2300) );
  OAI21X1 U27 ( .A(n1336), .B(n1330), .C(n2302), .Y(n3482) );
  NAND2X1 U28 ( .A(arr[5]), .B(n1337), .Y(n2302) );
  OAI21X1 U29 ( .A(n1336), .B(n1329), .C(n2304), .Y(n3483) );
  NAND2X1 U30 ( .A(arr[6]), .B(n1337), .Y(n2304) );
  OAI21X1 U31 ( .A(n1336), .B(n1328), .C(n2306), .Y(n3484) );
  NAND2X1 U32 ( .A(arr[7]), .B(n1337), .Y(n2306) );
  OAI21X1 U33 ( .A(n1336), .B(n1327), .C(n2308), .Y(n3485) );
  NAND2X1 U34 ( .A(arr[8]), .B(n1337), .Y(n2308) );
  OAI21X1 U35 ( .A(n1337), .B(n1326), .C(n2310), .Y(n3486) );
  NAND2X1 U36 ( .A(arr[9]), .B(n1337), .Y(n2310) );
  OAI21X1 U37 ( .A(n1337), .B(n1325), .C(n2312), .Y(n3487) );
  NAND2X1 U38 ( .A(arr[10]), .B(n1337), .Y(n2312) );
  OAI21X1 U39 ( .A(n1337), .B(n1324), .C(n2314), .Y(n3488) );
  NAND2X1 U40 ( .A(arr[11]), .B(n1337), .Y(n2314) );
  OAI21X1 U41 ( .A(n1336), .B(n1323), .C(n2316), .Y(n3489) );
  NAND2X1 U42 ( .A(arr[12]), .B(n1337), .Y(n2316) );
  OAI21X1 U43 ( .A(n1336), .B(n1322), .C(n2318), .Y(n3490) );
  NAND2X1 U44 ( .A(arr[13]), .B(n1337), .Y(n2318) );
  OAI21X1 U45 ( .A(n1336), .B(n1321), .C(n2320), .Y(n3491) );
  NAND2X1 U46 ( .A(arr[14]), .B(n1337), .Y(n2320) );
  OAI21X1 U47 ( .A(n1336), .B(n1320), .C(n2322), .Y(n3492) );
  NAND2X1 U48 ( .A(arr[15]), .B(n1337), .Y(n2322) );
  OAI21X1 U50 ( .A(n1335), .B(n1318), .C(n2326), .Y(n3493) );
  NAND2X1 U51 ( .A(arr[16]), .B(n1319), .Y(n2326) );
  OAI21X1 U52 ( .A(n1334), .B(n1318), .C(n2327), .Y(n3494) );
  NAND2X1 U53 ( .A(arr[17]), .B(n1319), .Y(n2327) );
  OAI21X1 U54 ( .A(n1333), .B(n1318), .C(n2328), .Y(n3495) );
  NAND2X1 U55 ( .A(arr[18]), .B(n1318), .Y(n2328) );
  OAI21X1 U56 ( .A(n1332), .B(n1318), .C(n2329), .Y(n3496) );
  NAND2X1 U57 ( .A(arr[19]), .B(n1318), .Y(n2329) );
  OAI21X1 U58 ( .A(n1331), .B(n1318), .C(n2330), .Y(n3497) );
  NAND2X1 U59 ( .A(arr[20]), .B(n1319), .Y(n2330) );
  OAI21X1 U60 ( .A(n1330), .B(n1318), .C(n2331), .Y(n3498) );
  NAND2X1 U61 ( .A(arr[21]), .B(n1319), .Y(n2331) );
  OAI21X1 U62 ( .A(n1329), .B(n1318), .C(n2332), .Y(n3499) );
  NAND2X1 U63 ( .A(arr[22]), .B(n1319), .Y(n2332) );
  OAI21X1 U64 ( .A(n1328), .B(n1318), .C(n2333), .Y(n3500) );
  NAND2X1 U65 ( .A(arr[23]), .B(n1319), .Y(n2333) );
  OAI21X1 U66 ( .A(n1327), .B(n1318), .C(n2334), .Y(n3501) );
  NAND2X1 U67 ( .A(arr[24]), .B(n1319), .Y(n2334) );
  OAI21X1 U68 ( .A(n1326), .B(n1319), .C(n2335), .Y(n3502) );
  NAND2X1 U69 ( .A(arr[25]), .B(n1319), .Y(n2335) );
  OAI21X1 U70 ( .A(n1325), .B(n1319), .C(n2336), .Y(n3503) );
  NAND2X1 U71 ( .A(arr[26]), .B(n1319), .Y(n2336) );
  OAI21X1 U72 ( .A(n1324), .B(n1319), .C(n2337), .Y(n3504) );
  NAND2X1 U73 ( .A(arr[27]), .B(n1319), .Y(n2337) );
  OAI21X1 U74 ( .A(n1323), .B(n1318), .C(n2338), .Y(n3505) );
  NAND2X1 U75 ( .A(arr[28]), .B(n1319), .Y(n2338) );
  OAI21X1 U76 ( .A(n1322), .B(n1318), .C(n2339), .Y(n3506) );
  NAND2X1 U77 ( .A(arr[29]), .B(n1319), .Y(n2339) );
  OAI21X1 U78 ( .A(n1321), .B(n1318), .C(n2340), .Y(n3507) );
  NAND2X1 U79 ( .A(arr[30]), .B(n1319), .Y(n2340) );
  OAI21X1 U80 ( .A(n1320), .B(n1318), .C(n2341), .Y(n3508) );
  NAND2X1 U81 ( .A(arr[31]), .B(n1319), .Y(n2341) );
  OAI21X1 U83 ( .A(n1335), .B(n1316), .C(n2344), .Y(n3509) );
  NAND2X1 U84 ( .A(arr[32]), .B(n1317), .Y(n2344) );
  OAI21X1 U85 ( .A(n1334), .B(n1316), .C(n2345), .Y(n3510) );
  NAND2X1 U86 ( .A(arr[33]), .B(n1317), .Y(n2345) );
  OAI21X1 U87 ( .A(n1333), .B(n1316), .C(n2346), .Y(n3511) );
  NAND2X1 U88 ( .A(arr[34]), .B(n1316), .Y(n2346) );
  OAI21X1 U89 ( .A(n1332), .B(n1316), .C(n2347), .Y(n3512) );
  NAND2X1 U90 ( .A(arr[35]), .B(n1316), .Y(n2347) );
  OAI21X1 U91 ( .A(n1331), .B(n1316), .C(n2348), .Y(n3513) );
  NAND2X1 U92 ( .A(arr[36]), .B(n1317), .Y(n2348) );
  OAI21X1 U93 ( .A(n1330), .B(n1316), .C(n2349), .Y(n3514) );
  NAND2X1 U94 ( .A(arr[37]), .B(n1317), .Y(n2349) );
  OAI21X1 U95 ( .A(n1329), .B(n1316), .C(n2350), .Y(n3515) );
  NAND2X1 U96 ( .A(arr[38]), .B(n1317), .Y(n2350) );
  OAI21X1 U97 ( .A(n1328), .B(n1316), .C(n2351), .Y(n3516) );
  NAND2X1 U98 ( .A(arr[39]), .B(n1317), .Y(n2351) );
  OAI21X1 U99 ( .A(n1327), .B(n1316), .C(n2352), .Y(n3517) );
  NAND2X1 U100 ( .A(arr[40]), .B(n1317), .Y(n2352) );
  OAI21X1 U101 ( .A(n1326), .B(n1317), .C(n2353), .Y(n3518) );
  NAND2X1 U102 ( .A(arr[41]), .B(n1317), .Y(n2353) );
  OAI21X1 U103 ( .A(n1325), .B(n1317), .C(n2354), .Y(n3519) );
  NAND2X1 U104 ( .A(arr[42]), .B(n1317), .Y(n2354) );
  OAI21X1 U105 ( .A(n1324), .B(n1317), .C(n2355), .Y(n3520) );
  NAND2X1 U106 ( .A(arr[43]), .B(n1317), .Y(n2355) );
  OAI21X1 U107 ( .A(n1323), .B(n1316), .C(n2356), .Y(n3521) );
  NAND2X1 U108 ( .A(arr[44]), .B(n1317), .Y(n2356) );
  OAI21X1 U109 ( .A(n1322), .B(n1316), .C(n2357), .Y(n3522) );
  NAND2X1 U110 ( .A(arr[45]), .B(n1317), .Y(n2357) );
  OAI21X1 U111 ( .A(n1321), .B(n1316), .C(n2358), .Y(n3523) );
  NAND2X1 U112 ( .A(arr[46]), .B(n1317), .Y(n2358) );
  OAI21X1 U113 ( .A(n1320), .B(n1316), .C(n2359), .Y(n3524) );
  NAND2X1 U114 ( .A(arr[47]), .B(n1317), .Y(n2359) );
  OAI21X1 U116 ( .A(n1335), .B(n1314), .C(n2362), .Y(n3525) );
  NAND2X1 U117 ( .A(arr[48]), .B(n1315), .Y(n2362) );
  OAI21X1 U118 ( .A(n1334), .B(n1314), .C(n2363), .Y(n3526) );
  NAND2X1 U119 ( .A(arr[49]), .B(n1315), .Y(n2363) );
  OAI21X1 U120 ( .A(n1333), .B(n1314), .C(n2364), .Y(n3527) );
  NAND2X1 U121 ( .A(arr[50]), .B(n1314), .Y(n2364) );
  OAI21X1 U122 ( .A(n1332), .B(n1314), .C(n2365), .Y(n3528) );
  NAND2X1 U123 ( .A(arr[51]), .B(n1314), .Y(n2365) );
  OAI21X1 U124 ( .A(n1331), .B(n1314), .C(n2366), .Y(n3529) );
  NAND2X1 U125 ( .A(arr[52]), .B(n1315), .Y(n2366) );
  OAI21X1 U126 ( .A(n1330), .B(n1314), .C(n2367), .Y(n3530) );
  NAND2X1 U127 ( .A(arr[53]), .B(n1315), .Y(n2367) );
  OAI21X1 U128 ( .A(n1329), .B(n1314), .C(n2368), .Y(n3531) );
  NAND2X1 U129 ( .A(arr[54]), .B(n1315), .Y(n2368) );
  OAI21X1 U130 ( .A(n1328), .B(n1314), .C(n2369), .Y(n3532) );
  NAND2X1 U131 ( .A(arr[55]), .B(n1315), .Y(n2369) );
  OAI21X1 U132 ( .A(n1327), .B(n1314), .C(n2370), .Y(n3533) );
  NAND2X1 U133 ( .A(arr[56]), .B(n1315), .Y(n2370) );
  OAI21X1 U134 ( .A(n1326), .B(n1315), .C(n2371), .Y(n3534) );
  NAND2X1 U135 ( .A(arr[57]), .B(n1315), .Y(n2371) );
  OAI21X1 U136 ( .A(n1325), .B(n1315), .C(n2372), .Y(n3535) );
  NAND2X1 U137 ( .A(arr[58]), .B(n1315), .Y(n2372) );
  OAI21X1 U138 ( .A(n1324), .B(n1315), .C(n2373), .Y(n3536) );
  NAND2X1 U139 ( .A(arr[59]), .B(n1315), .Y(n2373) );
  OAI21X1 U140 ( .A(n1323), .B(n1314), .C(n2374), .Y(n3537) );
  NAND2X1 U141 ( .A(arr[60]), .B(n1315), .Y(n2374) );
  OAI21X1 U142 ( .A(n1322), .B(n1314), .C(n2375), .Y(n3538) );
  NAND2X1 U143 ( .A(arr[61]), .B(n1315), .Y(n2375) );
  OAI21X1 U144 ( .A(n1321), .B(n1314), .C(n2376), .Y(n3539) );
  NAND2X1 U145 ( .A(arr[62]), .B(n1315), .Y(n2376) );
  OAI21X1 U146 ( .A(n1320), .B(n1314), .C(n2377), .Y(n3540) );
  NAND2X1 U147 ( .A(arr[63]), .B(n1315), .Y(n2377) );
  OAI21X1 U149 ( .A(n1335), .B(n1312), .C(n2379), .Y(n3541) );
  NAND2X1 U150 ( .A(arr[64]), .B(n1313), .Y(n2379) );
  OAI21X1 U151 ( .A(n1334), .B(n1312), .C(n2380), .Y(n3542) );
  NAND2X1 U152 ( .A(arr[65]), .B(n1313), .Y(n2380) );
  OAI21X1 U153 ( .A(n1333), .B(n1312), .C(n2381), .Y(n3543) );
  NAND2X1 U154 ( .A(arr[66]), .B(n1312), .Y(n2381) );
  OAI21X1 U155 ( .A(n1332), .B(n1312), .C(n2382), .Y(n3544) );
  NAND2X1 U156 ( .A(arr[67]), .B(n1312), .Y(n2382) );
  OAI21X1 U157 ( .A(n1331), .B(n1312), .C(n2383), .Y(n3545) );
  NAND2X1 U158 ( .A(arr[68]), .B(n1313), .Y(n2383) );
  OAI21X1 U159 ( .A(n1330), .B(n1312), .C(n2384), .Y(n3546) );
  NAND2X1 U160 ( .A(arr[69]), .B(n1313), .Y(n2384) );
  OAI21X1 U161 ( .A(n1329), .B(n1312), .C(n2385), .Y(n3547) );
  NAND2X1 U162 ( .A(arr[70]), .B(n1313), .Y(n2385) );
  OAI21X1 U163 ( .A(n1328), .B(n1312), .C(n2386), .Y(n3548) );
  NAND2X1 U164 ( .A(arr[71]), .B(n1313), .Y(n2386) );
  OAI21X1 U165 ( .A(n1327), .B(n1312), .C(n2387), .Y(n3549) );
  NAND2X1 U166 ( .A(arr[72]), .B(n1313), .Y(n2387) );
  OAI21X1 U167 ( .A(n1326), .B(n1313), .C(n2388), .Y(n3550) );
  NAND2X1 U168 ( .A(arr[73]), .B(n1313), .Y(n2388) );
  OAI21X1 U169 ( .A(n1325), .B(n1313), .C(n2389), .Y(n3551) );
  NAND2X1 U170 ( .A(arr[74]), .B(n1313), .Y(n2389) );
  OAI21X1 U171 ( .A(n1324), .B(n1313), .C(n2390), .Y(n3552) );
  NAND2X1 U172 ( .A(arr[75]), .B(n1313), .Y(n2390) );
  OAI21X1 U173 ( .A(n1323), .B(n1312), .C(n2391), .Y(n3553) );
  NAND2X1 U174 ( .A(arr[76]), .B(n1313), .Y(n2391) );
  OAI21X1 U175 ( .A(n1322), .B(n1312), .C(n2392), .Y(n3554) );
  NAND2X1 U176 ( .A(arr[77]), .B(n1313), .Y(n2392) );
  OAI21X1 U177 ( .A(n1321), .B(n1312), .C(n2393), .Y(n3555) );
  NAND2X1 U178 ( .A(arr[78]), .B(n1313), .Y(n2393) );
  OAI21X1 U179 ( .A(n1320), .B(n1312), .C(n2394), .Y(n3556) );
  NAND2X1 U180 ( .A(arr[79]), .B(n1313), .Y(n2394) );
  OAI21X1 U182 ( .A(n1335), .B(n1310), .C(n2397), .Y(n3557) );
  NAND2X1 U183 ( .A(arr[80]), .B(n1311), .Y(n2397) );
  OAI21X1 U184 ( .A(n1334), .B(n1310), .C(n2398), .Y(n3558) );
  NAND2X1 U185 ( .A(arr[81]), .B(n1311), .Y(n2398) );
  OAI21X1 U186 ( .A(n1333), .B(n1310), .C(n2399), .Y(n3559) );
  NAND2X1 U187 ( .A(arr[82]), .B(n1310), .Y(n2399) );
  OAI21X1 U188 ( .A(n1332), .B(n1310), .C(n2400), .Y(n3560) );
  NAND2X1 U189 ( .A(arr[83]), .B(n1310), .Y(n2400) );
  OAI21X1 U190 ( .A(n1331), .B(n1310), .C(n2401), .Y(n3561) );
  NAND2X1 U191 ( .A(arr[84]), .B(n1311), .Y(n2401) );
  OAI21X1 U192 ( .A(n1330), .B(n1310), .C(n2402), .Y(n3562) );
  NAND2X1 U193 ( .A(arr[85]), .B(n1311), .Y(n2402) );
  OAI21X1 U194 ( .A(n1329), .B(n1310), .C(n2403), .Y(n3563) );
  NAND2X1 U195 ( .A(arr[86]), .B(n1311), .Y(n2403) );
  OAI21X1 U196 ( .A(n1328), .B(n1310), .C(n2404), .Y(n3564) );
  NAND2X1 U197 ( .A(arr[87]), .B(n1311), .Y(n2404) );
  OAI21X1 U198 ( .A(n1327), .B(n1310), .C(n2405), .Y(n3565) );
  NAND2X1 U199 ( .A(arr[88]), .B(n1311), .Y(n2405) );
  OAI21X1 U200 ( .A(n1326), .B(n1311), .C(n2406), .Y(n3566) );
  NAND2X1 U201 ( .A(arr[89]), .B(n1311), .Y(n2406) );
  OAI21X1 U202 ( .A(n1325), .B(n1311), .C(n2407), .Y(n3567) );
  NAND2X1 U203 ( .A(arr[90]), .B(n1311), .Y(n2407) );
  OAI21X1 U204 ( .A(n1324), .B(n1311), .C(n2408), .Y(n3568) );
  NAND2X1 U205 ( .A(arr[91]), .B(n1311), .Y(n2408) );
  OAI21X1 U206 ( .A(n1323), .B(n1310), .C(n2409), .Y(n3569) );
  NAND2X1 U207 ( .A(arr[92]), .B(n1311), .Y(n2409) );
  OAI21X1 U208 ( .A(n1322), .B(n1310), .C(n2410), .Y(n3570) );
  NAND2X1 U209 ( .A(arr[93]), .B(n1311), .Y(n2410) );
  OAI21X1 U210 ( .A(n1321), .B(n1310), .C(n2411), .Y(n3571) );
  NAND2X1 U211 ( .A(arr[94]), .B(n1311), .Y(n2411) );
  OAI21X1 U212 ( .A(n1320), .B(n1310), .C(n2412), .Y(n3572) );
  NAND2X1 U213 ( .A(arr[95]), .B(n1311), .Y(n2412) );
  OAI21X1 U215 ( .A(n1335), .B(n1308), .C(n2414), .Y(n3573) );
  NAND2X1 U216 ( .A(arr[96]), .B(n1309), .Y(n2414) );
  OAI21X1 U217 ( .A(n1334), .B(n1308), .C(n2415), .Y(n3574) );
  NAND2X1 U218 ( .A(arr[97]), .B(n1309), .Y(n2415) );
  OAI21X1 U219 ( .A(n1333), .B(n1308), .C(n2416), .Y(n3575) );
  NAND2X1 U220 ( .A(arr[98]), .B(n1308), .Y(n2416) );
  OAI21X1 U221 ( .A(n1332), .B(n1308), .C(n2417), .Y(n3576) );
  NAND2X1 U222 ( .A(arr[99]), .B(n1308), .Y(n2417) );
  OAI21X1 U223 ( .A(n1331), .B(n1308), .C(n2418), .Y(n3577) );
  NAND2X1 U224 ( .A(arr[100]), .B(n1309), .Y(n2418) );
  OAI21X1 U225 ( .A(n1330), .B(n1308), .C(n2419), .Y(n3578) );
  NAND2X1 U226 ( .A(arr[101]), .B(n1309), .Y(n2419) );
  OAI21X1 U227 ( .A(n1329), .B(n1308), .C(n2420), .Y(n3579) );
  NAND2X1 U228 ( .A(arr[102]), .B(n1309), .Y(n2420) );
  OAI21X1 U229 ( .A(n1328), .B(n1308), .C(n2421), .Y(n3580) );
  NAND2X1 U230 ( .A(arr[103]), .B(n1309), .Y(n2421) );
  OAI21X1 U231 ( .A(n1327), .B(n1308), .C(n2422), .Y(n3581) );
  NAND2X1 U232 ( .A(arr[104]), .B(n1309), .Y(n2422) );
  OAI21X1 U233 ( .A(n1326), .B(n1309), .C(n2423), .Y(n3582) );
  NAND2X1 U234 ( .A(arr[105]), .B(n1309), .Y(n2423) );
  OAI21X1 U235 ( .A(n1325), .B(n1309), .C(n2424), .Y(n3583) );
  NAND2X1 U236 ( .A(arr[106]), .B(n1309), .Y(n2424) );
  OAI21X1 U237 ( .A(n1324), .B(n1309), .C(n2425), .Y(n3584) );
  NAND2X1 U238 ( .A(arr[107]), .B(n1309), .Y(n2425) );
  OAI21X1 U239 ( .A(n1323), .B(n1308), .C(n2426), .Y(n3585) );
  NAND2X1 U240 ( .A(arr[108]), .B(n1309), .Y(n2426) );
  OAI21X1 U241 ( .A(n1322), .B(n1308), .C(n2427), .Y(n3586) );
  NAND2X1 U242 ( .A(arr[109]), .B(n1309), .Y(n2427) );
  OAI21X1 U243 ( .A(n1321), .B(n1308), .C(n2428), .Y(n3587) );
  NAND2X1 U244 ( .A(arr[110]), .B(n1309), .Y(n2428) );
  OAI21X1 U245 ( .A(n1320), .B(n1308), .C(n2429), .Y(n3588) );
  NAND2X1 U246 ( .A(arr[111]), .B(n1309), .Y(n2429) );
  OAI21X1 U248 ( .A(n1335), .B(n1306), .C(n2432), .Y(n3589) );
  NAND2X1 U249 ( .A(arr[112]), .B(n1307), .Y(n2432) );
  OAI21X1 U250 ( .A(n1334), .B(n1306), .C(n2433), .Y(n3590) );
  NAND2X1 U251 ( .A(arr[113]), .B(n1307), .Y(n2433) );
  OAI21X1 U252 ( .A(n1333), .B(n1306), .C(n2434), .Y(n3591) );
  NAND2X1 U253 ( .A(arr[114]), .B(n1306), .Y(n2434) );
  OAI21X1 U254 ( .A(n1332), .B(n1306), .C(n2435), .Y(n3592) );
  NAND2X1 U255 ( .A(arr[115]), .B(n1306), .Y(n2435) );
  OAI21X1 U256 ( .A(n1331), .B(n1306), .C(n2436), .Y(n3593) );
  NAND2X1 U257 ( .A(arr[116]), .B(n1307), .Y(n2436) );
  OAI21X1 U258 ( .A(n1330), .B(n1306), .C(n2437), .Y(n3594) );
  NAND2X1 U259 ( .A(arr[117]), .B(n1307), .Y(n2437) );
  OAI21X1 U260 ( .A(n1329), .B(n1306), .C(n2438), .Y(n3595) );
  NAND2X1 U261 ( .A(arr[118]), .B(n1307), .Y(n2438) );
  OAI21X1 U262 ( .A(n1328), .B(n1306), .C(n2439), .Y(n3596) );
  NAND2X1 U263 ( .A(arr[119]), .B(n1307), .Y(n2439) );
  OAI21X1 U264 ( .A(n1327), .B(n1306), .C(n2440), .Y(n3597) );
  NAND2X1 U265 ( .A(arr[120]), .B(n1307), .Y(n2440) );
  OAI21X1 U266 ( .A(n1326), .B(n1307), .C(n2441), .Y(n3598) );
  NAND2X1 U267 ( .A(arr[121]), .B(n1307), .Y(n2441) );
  OAI21X1 U268 ( .A(n1325), .B(n1307), .C(n2442), .Y(n3599) );
  NAND2X1 U269 ( .A(arr[122]), .B(n1307), .Y(n2442) );
  OAI21X1 U270 ( .A(n1324), .B(n1307), .C(n2443), .Y(n3600) );
  NAND2X1 U271 ( .A(arr[123]), .B(n1307), .Y(n2443) );
  OAI21X1 U272 ( .A(n1323), .B(n1306), .C(n2444), .Y(n3601) );
  NAND2X1 U273 ( .A(arr[124]), .B(n1307), .Y(n2444) );
  OAI21X1 U274 ( .A(n1322), .B(n1306), .C(n2445), .Y(n3602) );
  NAND2X1 U275 ( .A(arr[125]), .B(n1307), .Y(n2445) );
  OAI21X1 U276 ( .A(n1321), .B(n1306), .C(n2446), .Y(n3603) );
  NAND2X1 U277 ( .A(arr[126]), .B(n1307), .Y(n2446) );
  OAI21X1 U278 ( .A(n1320), .B(n1306), .C(n2447), .Y(n3604) );
  NAND2X1 U279 ( .A(arr[127]), .B(n1307), .Y(n2447) );
  OAI21X1 U281 ( .A(n1335), .B(n1304), .C(n2449), .Y(n3605) );
  NAND2X1 U282 ( .A(arr[128]), .B(n1305), .Y(n2449) );
  OAI21X1 U283 ( .A(n1334), .B(n1304), .C(n2450), .Y(n3606) );
  NAND2X1 U284 ( .A(arr[129]), .B(n1305), .Y(n2450) );
  OAI21X1 U285 ( .A(n1333), .B(n1304), .C(n2451), .Y(n3607) );
  NAND2X1 U286 ( .A(arr[130]), .B(n1304), .Y(n2451) );
  OAI21X1 U287 ( .A(n1332), .B(n1304), .C(n2452), .Y(n3608) );
  NAND2X1 U288 ( .A(arr[131]), .B(n1304), .Y(n2452) );
  OAI21X1 U289 ( .A(n1331), .B(n1304), .C(n2453), .Y(n3609) );
  NAND2X1 U290 ( .A(arr[132]), .B(n1305), .Y(n2453) );
  OAI21X1 U291 ( .A(n1330), .B(n1304), .C(n2454), .Y(n3610) );
  NAND2X1 U292 ( .A(arr[133]), .B(n1305), .Y(n2454) );
  OAI21X1 U293 ( .A(n1329), .B(n1304), .C(n2455), .Y(n3611) );
  NAND2X1 U294 ( .A(arr[134]), .B(n1305), .Y(n2455) );
  OAI21X1 U295 ( .A(n1328), .B(n1304), .C(n2456), .Y(n3612) );
  NAND2X1 U296 ( .A(arr[135]), .B(n1305), .Y(n2456) );
  OAI21X1 U297 ( .A(n1327), .B(n1304), .C(n2457), .Y(n3613) );
  NAND2X1 U298 ( .A(arr[136]), .B(n1305), .Y(n2457) );
  OAI21X1 U299 ( .A(n1326), .B(n1305), .C(n2458), .Y(n3614) );
  NAND2X1 U300 ( .A(arr[137]), .B(n1305), .Y(n2458) );
  OAI21X1 U301 ( .A(n1325), .B(n1305), .C(n2459), .Y(n3615) );
  NAND2X1 U302 ( .A(arr[138]), .B(n1305), .Y(n2459) );
  OAI21X1 U303 ( .A(n1324), .B(n1305), .C(n2460), .Y(n3616) );
  NAND2X1 U304 ( .A(arr[139]), .B(n1305), .Y(n2460) );
  OAI21X1 U305 ( .A(n1323), .B(n1304), .C(n2461), .Y(n3617) );
  NAND2X1 U306 ( .A(arr[140]), .B(n1305), .Y(n2461) );
  OAI21X1 U307 ( .A(n1322), .B(n1304), .C(n2462), .Y(n3618) );
  NAND2X1 U308 ( .A(arr[141]), .B(n1305), .Y(n2462) );
  OAI21X1 U309 ( .A(n1321), .B(n1304), .C(n2463), .Y(n3619) );
  NAND2X1 U310 ( .A(arr[142]), .B(n1305), .Y(n2463) );
  OAI21X1 U311 ( .A(n1320), .B(n1304), .C(n2464), .Y(n3620) );
  NAND2X1 U312 ( .A(arr[143]), .B(n1305), .Y(n2464) );
  OAI21X1 U314 ( .A(n1335), .B(n1302), .C(n2467), .Y(n3621) );
  NAND2X1 U315 ( .A(arr[144]), .B(n1303), .Y(n2467) );
  OAI21X1 U316 ( .A(n1334), .B(n1302), .C(n2468), .Y(n3622) );
  NAND2X1 U317 ( .A(arr[145]), .B(n1303), .Y(n2468) );
  OAI21X1 U318 ( .A(n1333), .B(n1302), .C(n2469), .Y(n3623) );
  NAND2X1 U319 ( .A(arr[146]), .B(n1302), .Y(n2469) );
  OAI21X1 U320 ( .A(n1332), .B(n1302), .C(n2470), .Y(n3624) );
  NAND2X1 U321 ( .A(arr[147]), .B(n1302), .Y(n2470) );
  OAI21X1 U322 ( .A(n1331), .B(n1302), .C(n2471), .Y(n3625) );
  NAND2X1 U323 ( .A(arr[148]), .B(n1303), .Y(n2471) );
  OAI21X1 U324 ( .A(n1330), .B(n1302), .C(n2472), .Y(n3626) );
  NAND2X1 U325 ( .A(arr[149]), .B(n1303), .Y(n2472) );
  OAI21X1 U326 ( .A(n1329), .B(n1302), .C(n2473), .Y(n3627) );
  NAND2X1 U327 ( .A(arr[150]), .B(n1303), .Y(n2473) );
  OAI21X1 U328 ( .A(n1328), .B(n1302), .C(n2474), .Y(n3628) );
  NAND2X1 U329 ( .A(arr[151]), .B(n1303), .Y(n2474) );
  OAI21X1 U330 ( .A(n1327), .B(n1302), .C(n2475), .Y(n3629) );
  NAND2X1 U331 ( .A(arr[152]), .B(n1303), .Y(n2475) );
  OAI21X1 U332 ( .A(n1326), .B(n1303), .C(n2476), .Y(n3630) );
  NAND2X1 U333 ( .A(arr[153]), .B(n1303), .Y(n2476) );
  OAI21X1 U334 ( .A(n1325), .B(n1303), .C(n2477), .Y(n3631) );
  NAND2X1 U335 ( .A(arr[154]), .B(n1303), .Y(n2477) );
  OAI21X1 U336 ( .A(n1324), .B(n1303), .C(n2478), .Y(n3632) );
  NAND2X1 U337 ( .A(arr[155]), .B(n1303), .Y(n2478) );
  OAI21X1 U338 ( .A(n1323), .B(n1302), .C(n2479), .Y(n3633) );
  NAND2X1 U339 ( .A(arr[156]), .B(n1303), .Y(n2479) );
  OAI21X1 U340 ( .A(n1322), .B(n1302), .C(n2480), .Y(n3634) );
  NAND2X1 U341 ( .A(arr[157]), .B(n1303), .Y(n2480) );
  OAI21X1 U342 ( .A(n1321), .B(n1302), .C(n2481), .Y(n3635) );
  NAND2X1 U343 ( .A(arr[158]), .B(n1303), .Y(n2481) );
  OAI21X1 U344 ( .A(n1320), .B(n1302), .C(n2482), .Y(n3636) );
  NAND2X1 U345 ( .A(arr[159]), .B(n1303), .Y(n2482) );
  OAI21X1 U347 ( .A(n1335), .B(n1300), .C(n2484), .Y(n3637) );
  NAND2X1 U348 ( .A(arr[160]), .B(n1301), .Y(n2484) );
  OAI21X1 U349 ( .A(n1334), .B(n1300), .C(n2485), .Y(n3638) );
  NAND2X1 U350 ( .A(arr[161]), .B(n1301), .Y(n2485) );
  OAI21X1 U351 ( .A(n1333), .B(n1300), .C(n2486), .Y(n3639) );
  NAND2X1 U352 ( .A(arr[162]), .B(n1300), .Y(n2486) );
  OAI21X1 U353 ( .A(n1332), .B(n1300), .C(n2487), .Y(n3640) );
  NAND2X1 U354 ( .A(arr[163]), .B(n1300), .Y(n2487) );
  OAI21X1 U355 ( .A(n1331), .B(n1300), .C(n2488), .Y(n3641) );
  NAND2X1 U356 ( .A(arr[164]), .B(n1301), .Y(n2488) );
  OAI21X1 U357 ( .A(n1330), .B(n1300), .C(n2489), .Y(n3642) );
  NAND2X1 U358 ( .A(arr[165]), .B(n1301), .Y(n2489) );
  OAI21X1 U359 ( .A(n1329), .B(n1300), .C(n2490), .Y(n3643) );
  NAND2X1 U360 ( .A(arr[166]), .B(n1301), .Y(n2490) );
  OAI21X1 U361 ( .A(n1328), .B(n1300), .C(n2491), .Y(n3644) );
  NAND2X1 U362 ( .A(arr[167]), .B(n1301), .Y(n2491) );
  OAI21X1 U363 ( .A(n1327), .B(n1300), .C(n2492), .Y(n3645) );
  NAND2X1 U364 ( .A(arr[168]), .B(n1301), .Y(n2492) );
  OAI21X1 U365 ( .A(n1326), .B(n1301), .C(n2493), .Y(n3646) );
  NAND2X1 U366 ( .A(arr[169]), .B(n1301), .Y(n2493) );
  OAI21X1 U367 ( .A(n1325), .B(n1301), .C(n2494), .Y(n3647) );
  NAND2X1 U368 ( .A(arr[170]), .B(n1301), .Y(n2494) );
  OAI21X1 U369 ( .A(n1324), .B(n1301), .C(n2495), .Y(n3648) );
  NAND2X1 U370 ( .A(arr[171]), .B(n1301), .Y(n2495) );
  OAI21X1 U371 ( .A(n1323), .B(n1300), .C(n2496), .Y(n3649) );
  NAND2X1 U372 ( .A(arr[172]), .B(n1301), .Y(n2496) );
  OAI21X1 U373 ( .A(n1322), .B(n1300), .C(n2497), .Y(n3650) );
  NAND2X1 U374 ( .A(arr[173]), .B(n1301), .Y(n2497) );
  OAI21X1 U375 ( .A(n1321), .B(n1300), .C(n2498), .Y(n3651) );
  NAND2X1 U376 ( .A(arr[174]), .B(n1301), .Y(n2498) );
  OAI21X1 U377 ( .A(n1320), .B(n1300), .C(n2499), .Y(n3652) );
  NAND2X1 U378 ( .A(arr[175]), .B(n1301), .Y(n2499) );
  OAI21X1 U380 ( .A(n1335), .B(n1298), .C(n2502), .Y(n3653) );
  NAND2X1 U381 ( .A(arr[176]), .B(n1299), .Y(n2502) );
  OAI21X1 U382 ( .A(n1334), .B(n1298), .C(n2503), .Y(n3654) );
  NAND2X1 U383 ( .A(arr[177]), .B(n1299), .Y(n2503) );
  OAI21X1 U384 ( .A(n1333), .B(n1298), .C(n2504), .Y(n3655) );
  NAND2X1 U385 ( .A(arr[178]), .B(n1298), .Y(n2504) );
  OAI21X1 U386 ( .A(n1332), .B(n1298), .C(n2505), .Y(n3656) );
  NAND2X1 U387 ( .A(arr[179]), .B(n1298), .Y(n2505) );
  OAI21X1 U388 ( .A(n1331), .B(n1298), .C(n2506), .Y(n3657) );
  NAND2X1 U389 ( .A(arr[180]), .B(n1299), .Y(n2506) );
  OAI21X1 U390 ( .A(n1330), .B(n1298), .C(n2507), .Y(n3658) );
  NAND2X1 U391 ( .A(arr[181]), .B(n1299), .Y(n2507) );
  OAI21X1 U392 ( .A(n1329), .B(n1298), .C(n2508), .Y(n3659) );
  NAND2X1 U393 ( .A(arr[182]), .B(n1299), .Y(n2508) );
  OAI21X1 U394 ( .A(n1328), .B(n1298), .C(n2509), .Y(n3660) );
  NAND2X1 U395 ( .A(arr[183]), .B(n1299), .Y(n2509) );
  OAI21X1 U396 ( .A(n1327), .B(n1298), .C(n2510), .Y(n3661) );
  NAND2X1 U397 ( .A(arr[184]), .B(n1299), .Y(n2510) );
  OAI21X1 U398 ( .A(n1326), .B(n1299), .C(n2511), .Y(n3662) );
  NAND2X1 U399 ( .A(arr[185]), .B(n1299), .Y(n2511) );
  OAI21X1 U400 ( .A(n1325), .B(n1299), .C(n2512), .Y(n3663) );
  NAND2X1 U401 ( .A(arr[186]), .B(n1299), .Y(n2512) );
  OAI21X1 U402 ( .A(n1324), .B(n1299), .C(n2513), .Y(n3664) );
  NAND2X1 U403 ( .A(arr[187]), .B(n1299), .Y(n2513) );
  OAI21X1 U404 ( .A(n1323), .B(n1298), .C(n2514), .Y(n3665) );
  NAND2X1 U405 ( .A(arr[188]), .B(n1299), .Y(n2514) );
  OAI21X1 U406 ( .A(n1322), .B(n1298), .C(n2515), .Y(n3666) );
  NAND2X1 U407 ( .A(arr[189]), .B(n1299), .Y(n2515) );
  OAI21X1 U408 ( .A(n1321), .B(n1298), .C(n2516), .Y(n3667) );
  NAND2X1 U409 ( .A(arr[190]), .B(n1299), .Y(n2516) );
  OAI21X1 U410 ( .A(n1320), .B(n1298), .C(n2517), .Y(n3668) );
  NAND2X1 U411 ( .A(arr[191]), .B(n1299), .Y(n2517) );
  OAI21X1 U413 ( .A(n1335), .B(n1296), .C(n2519), .Y(n3669) );
  NAND2X1 U414 ( .A(arr[192]), .B(n1297), .Y(n2519) );
  OAI21X1 U415 ( .A(n1334), .B(n1296), .C(n2520), .Y(n3670) );
  NAND2X1 U416 ( .A(arr[193]), .B(n1297), .Y(n2520) );
  OAI21X1 U417 ( .A(n1333), .B(n1296), .C(n2521), .Y(n3671) );
  NAND2X1 U418 ( .A(arr[194]), .B(n1296), .Y(n2521) );
  OAI21X1 U419 ( .A(n1332), .B(n1296), .C(n2522), .Y(n3672) );
  NAND2X1 U420 ( .A(arr[195]), .B(n1296), .Y(n2522) );
  OAI21X1 U421 ( .A(n1331), .B(n1296), .C(n2523), .Y(n3673) );
  NAND2X1 U422 ( .A(arr[196]), .B(n1297), .Y(n2523) );
  OAI21X1 U423 ( .A(n1330), .B(n1296), .C(n2524), .Y(n3674) );
  NAND2X1 U424 ( .A(arr[197]), .B(n1297), .Y(n2524) );
  OAI21X1 U425 ( .A(n1329), .B(n1296), .C(n2525), .Y(n3675) );
  NAND2X1 U426 ( .A(arr[198]), .B(n1297), .Y(n2525) );
  OAI21X1 U427 ( .A(n1328), .B(n1296), .C(n2526), .Y(n3676) );
  NAND2X1 U428 ( .A(arr[199]), .B(n1297), .Y(n2526) );
  OAI21X1 U429 ( .A(n1327), .B(n1296), .C(n2527), .Y(n3677) );
  NAND2X1 U430 ( .A(arr[200]), .B(n1297), .Y(n2527) );
  OAI21X1 U431 ( .A(n1326), .B(n1297), .C(n2528), .Y(n3678) );
  NAND2X1 U432 ( .A(arr[201]), .B(n1297), .Y(n2528) );
  OAI21X1 U433 ( .A(n1325), .B(n1297), .C(n2529), .Y(n3679) );
  NAND2X1 U434 ( .A(arr[202]), .B(n1297), .Y(n2529) );
  OAI21X1 U435 ( .A(n1324), .B(n1297), .C(n2530), .Y(n3680) );
  NAND2X1 U436 ( .A(arr[203]), .B(n1297), .Y(n2530) );
  OAI21X1 U437 ( .A(n1323), .B(n1296), .C(n2531), .Y(n3681) );
  NAND2X1 U438 ( .A(arr[204]), .B(n1297), .Y(n2531) );
  OAI21X1 U439 ( .A(n1322), .B(n1296), .C(n2532), .Y(n3682) );
  NAND2X1 U440 ( .A(arr[205]), .B(n1297), .Y(n2532) );
  OAI21X1 U441 ( .A(n1321), .B(n1296), .C(n2533), .Y(n3683) );
  NAND2X1 U442 ( .A(arr[206]), .B(n1297), .Y(n2533) );
  OAI21X1 U443 ( .A(n1320), .B(n1296), .C(n2534), .Y(n3684) );
  NAND2X1 U444 ( .A(arr[207]), .B(n1297), .Y(n2534) );
  OAI21X1 U446 ( .A(n1335), .B(n1294), .C(n2537), .Y(n3685) );
  NAND2X1 U447 ( .A(arr[208]), .B(n1295), .Y(n2537) );
  OAI21X1 U448 ( .A(n1334), .B(n1294), .C(n2538), .Y(n3686) );
  NAND2X1 U449 ( .A(arr[209]), .B(n1295), .Y(n2538) );
  OAI21X1 U450 ( .A(n1333), .B(n1294), .C(n2539), .Y(n3687) );
  NAND2X1 U451 ( .A(arr[210]), .B(n1294), .Y(n2539) );
  OAI21X1 U452 ( .A(n1332), .B(n1294), .C(n2540), .Y(n3688) );
  NAND2X1 U453 ( .A(arr[211]), .B(n1294), .Y(n2540) );
  OAI21X1 U454 ( .A(n1331), .B(n1294), .C(n2541), .Y(n3689) );
  NAND2X1 U455 ( .A(arr[212]), .B(n1295), .Y(n2541) );
  OAI21X1 U456 ( .A(n1330), .B(n1294), .C(n2542), .Y(n3690) );
  NAND2X1 U457 ( .A(arr[213]), .B(n1295), .Y(n2542) );
  OAI21X1 U458 ( .A(n1329), .B(n1294), .C(n2543), .Y(n3691) );
  NAND2X1 U459 ( .A(arr[214]), .B(n1295), .Y(n2543) );
  OAI21X1 U460 ( .A(n1328), .B(n1294), .C(n2544), .Y(n3692) );
  NAND2X1 U461 ( .A(arr[215]), .B(n1295), .Y(n2544) );
  OAI21X1 U462 ( .A(n1327), .B(n1294), .C(n2545), .Y(n3693) );
  NAND2X1 U463 ( .A(arr[216]), .B(n1295), .Y(n2545) );
  OAI21X1 U464 ( .A(n1326), .B(n1295), .C(n2546), .Y(n3694) );
  NAND2X1 U465 ( .A(arr[217]), .B(n1295), .Y(n2546) );
  OAI21X1 U466 ( .A(n1325), .B(n1295), .C(n2547), .Y(n3695) );
  NAND2X1 U467 ( .A(arr[218]), .B(n1295), .Y(n2547) );
  OAI21X1 U468 ( .A(n1324), .B(n1295), .C(n2548), .Y(n3696) );
  NAND2X1 U469 ( .A(arr[219]), .B(n1295), .Y(n2548) );
  OAI21X1 U470 ( .A(n1323), .B(n1294), .C(n2549), .Y(n3697) );
  NAND2X1 U471 ( .A(arr[220]), .B(n1295), .Y(n2549) );
  OAI21X1 U472 ( .A(n1322), .B(n1294), .C(n2550), .Y(n3698) );
  NAND2X1 U473 ( .A(arr[221]), .B(n1295), .Y(n2550) );
  OAI21X1 U474 ( .A(n1321), .B(n1294), .C(n2551), .Y(n3699) );
  NAND2X1 U475 ( .A(arr[222]), .B(n1295), .Y(n2551) );
  OAI21X1 U476 ( .A(n1320), .B(n1294), .C(n2552), .Y(n3700) );
  NAND2X1 U477 ( .A(arr[223]), .B(n1295), .Y(n2552) );
  OAI21X1 U479 ( .A(n1335), .B(n1292), .C(n2554), .Y(n3701) );
  NAND2X1 U480 ( .A(arr[224]), .B(n1293), .Y(n2554) );
  OAI21X1 U481 ( .A(n1334), .B(n1292), .C(n2555), .Y(n3702) );
  NAND2X1 U482 ( .A(arr[225]), .B(n1293), .Y(n2555) );
  OAI21X1 U483 ( .A(n1333), .B(n1292), .C(n2556), .Y(n3703) );
  NAND2X1 U484 ( .A(arr[226]), .B(n1292), .Y(n2556) );
  OAI21X1 U485 ( .A(n1332), .B(n1292), .C(n2557), .Y(n3704) );
  NAND2X1 U486 ( .A(arr[227]), .B(n1292), .Y(n2557) );
  OAI21X1 U487 ( .A(n1331), .B(n1292), .C(n2558), .Y(n3705) );
  NAND2X1 U488 ( .A(arr[228]), .B(n1293), .Y(n2558) );
  OAI21X1 U489 ( .A(n1330), .B(n1292), .C(n2559), .Y(n3706) );
  NAND2X1 U490 ( .A(arr[229]), .B(n1293), .Y(n2559) );
  OAI21X1 U491 ( .A(n1329), .B(n1292), .C(n2560), .Y(n3707) );
  NAND2X1 U492 ( .A(arr[230]), .B(n1293), .Y(n2560) );
  OAI21X1 U493 ( .A(n1328), .B(n1292), .C(n2561), .Y(n3708) );
  NAND2X1 U494 ( .A(arr[231]), .B(n1293), .Y(n2561) );
  OAI21X1 U495 ( .A(n1327), .B(n1292), .C(n2562), .Y(n3709) );
  NAND2X1 U496 ( .A(arr[232]), .B(n1293), .Y(n2562) );
  OAI21X1 U497 ( .A(n1326), .B(n1293), .C(n2563), .Y(n3710) );
  NAND2X1 U498 ( .A(arr[233]), .B(n1293), .Y(n2563) );
  OAI21X1 U499 ( .A(n1325), .B(n1293), .C(n2564), .Y(n3711) );
  NAND2X1 U500 ( .A(arr[234]), .B(n1293), .Y(n2564) );
  OAI21X1 U501 ( .A(n1324), .B(n1293), .C(n2565), .Y(n3712) );
  NAND2X1 U502 ( .A(arr[235]), .B(n1293), .Y(n2565) );
  OAI21X1 U503 ( .A(n1323), .B(n1292), .C(n2566), .Y(n3713) );
  NAND2X1 U504 ( .A(arr[236]), .B(n1293), .Y(n2566) );
  OAI21X1 U505 ( .A(n1322), .B(n1292), .C(n2567), .Y(n3714) );
  NAND2X1 U506 ( .A(arr[237]), .B(n1293), .Y(n2567) );
  OAI21X1 U507 ( .A(n1321), .B(n1292), .C(n2568), .Y(n3715) );
  NAND2X1 U508 ( .A(arr[238]), .B(n1293), .Y(n2568) );
  OAI21X1 U509 ( .A(n1320), .B(n1292), .C(n2569), .Y(n3716) );
  NAND2X1 U510 ( .A(arr[239]), .B(n1293), .Y(n2569) );
  OAI21X1 U512 ( .A(n1335), .B(n1290), .C(n2572), .Y(n3717) );
  NAND2X1 U513 ( .A(arr[240]), .B(n1291), .Y(n2572) );
  OAI21X1 U514 ( .A(n1334), .B(n1290), .C(n2573), .Y(n3718) );
  NAND2X1 U515 ( .A(arr[241]), .B(n1291), .Y(n2573) );
  OAI21X1 U516 ( .A(n1333), .B(n1290), .C(n2574), .Y(n3719) );
  NAND2X1 U517 ( .A(arr[242]), .B(n1290), .Y(n2574) );
  OAI21X1 U518 ( .A(n1332), .B(n1290), .C(n2575), .Y(n3720) );
  NAND2X1 U519 ( .A(arr[243]), .B(n1290), .Y(n2575) );
  OAI21X1 U520 ( .A(n1331), .B(n1290), .C(n2576), .Y(n3721) );
  NAND2X1 U521 ( .A(arr[244]), .B(n1291), .Y(n2576) );
  OAI21X1 U522 ( .A(n1330), .B(n1290), .C(n2577), .Y(n3722) );
  NAND2X1 U523 ( .A(arr[245]), .B(n1291), .Y(n2577) );
  OAI21X1 U524 ( .A(n1329), .B(n1290), .C(n2578), .Y(n3723) );
  NAND2X1 U525 ( .A(arr[246]), .B(n1291), .Y(n2578) );
  OAI21X1 U526 ( .A(n1328), .B(n1290), .C(n2579), .Y(n3724) );
  NAND2X1 U527 ( .A(arr[247]), .B(n1291), .Y(n2579) );
  OAI21X1 U528 ( .A(n1327), .B(n1290), .C(n2580), .Y(n3725) );
  NAND2X1 U529 ( .A(arr[248]), .B(n1291), .Y(n2580) );
  OAI21X1 U530 ( .A(n1326), .B(n1291), .C(n2581), .Y(n3726) );
  NAND2X1 U531 ( .A(arr[249]), .B(n1291), .Y(n2581) );
  OAI21X1 U532 ( .A(n1325), .B(n1291), .C(n2582), .Y(n3727) );
  NAND2X1 U533 ( .A(arr[250]), .B(n1291), .Y(n2582) );
  OAI21X1 U534 ( .A(n1324), .B(n1291), .C(n2583), .Y(n3728) );
  NAND2X1 U535 ( .A(arr[251]), .B(n1291), .Y(n2583) );
  OAI21X1 U536 ( .A(n1323), .B(n1290), .C(n2584), .Y(n3729) );
  NAND2X1 U537 ( .A(arr[252]), .B(n1291), .Y(n2584) );
  OAI21X1 U538 ( .A(n1322), .B(n1290), .C(n2585), .Y(n3730) );
  NAND2X1 U539 ( .A(arr[253]), .B(n1291), .Y(n2585) );
  OAI21X1 U540 ( .A(n1321), .B(n1290), .C(n2586), .Y(n3731) );
  NAND2X1 U541 ( .A(arr[254]), .B(n1291), .Y(n2586) );
  OAI21X1 U542 ( .A(n1320), .B(n1290), .C(n2587), .Y(n3732) );
  NAND2X1 U543 ( .A(arr[255]), .B(n1291), .Y(n2587) );
  OAI21X1 U545 ( .A(n1335), .B(n1288), .C(n2589), .Y(n3733) );
  NAND2X1 U546 ( .A(arr[256]), .B(n1289), .Y(n2589) );
  OAI21X1 U547 ( .A(n1334), .B(n1288), .C(n2590), .Y(n3734) );
  NAND2X1 U548 ( .A(arr[257]), .B(n1289), .Y(n2590) );
  OAI21X1 U549 ( .A(n1333), .B(n1288), .C(n2591), .Y(n3735) );
  NAND2X1 U550 ( .A(arr[258]), .B(n1288), .Y(n2591) );
  OAI21X1 U551 ( .A(n1332), .B(n1288), .C(n2592), .Y(n3736) );
  NAND2X1 U552 ( .A(arr[259]), .B(n1288), .Y(n2592) );
  OAI21X1 U553 ( .A(n1331), .B(n1288), .C(n2593), .Y(n3737) );
  NAND2X1 U554 ( .A(arr[260]), .B(n1289), .Y(n2593) );
  OAI21X1 U555 ( .A(n1330), .B(n1288), .C(n2594), .Y(n3738) );
  NAND2X1 U556 ( .A(arr[261]), .B(n1289), .Y(n2594) );
  OAI21X1 U557 ( .A(n1329), .B(n1288), .C(n2595), .Y(n3739) );
  NAND2X1 U558 ( .A(arr[262]), .B(n1289), .Y(n2595) );
  OAI21X1 U559 ( .A(n1328), .B(n1288), .C(n2596), .Y(n3740) );
  NAND2X1 U560 ( .A(arr[263]), .B(n1289), .Y(n2596) );
  OAI21X1 U561 ( .A(n1327), .B(n1288), .C(n2597), .Y(n3741) );
  NAND2X1 U562 ( .A(arr[264]), .B(n1289), .Y(n2597) );
  OAI21X1 U563 ( .A(n1326), .B(n1289), .C(n2598), .Y(n3742) );
  NAND2X1 U564 ( .A(arr[265]), .B(n1289), .Y(n2598) );
  OAI21X1 U565 ( .A(n1325), .B(n1289), .C(n2599), .Y(n3743) );
  NAND2X1 U566 ( .A(arr[266]), .B(n1289), .Y(n2599) );
  OAI21X1 U567 ( .A(n1324), .B(n1289), .C(n2600), .Y(n3744) );
  NAND2X1 U568 ( .A(arr[267]), .B(n1289), .Y(n2600) );
  OAI21X1 U569 ( .A(n1323), .B(n1288), .C(n2601), .Y(n3745) );
  NAND2X1 U570 ( .A(arr[268]), .B(n1289), .Y(n2601) );
  OAI21X1 U571 ( .A(n1322), .B(n1288), .C(n2602), .Y(n3746) );
  NAND2X1 U572 ( .A(arr[269]), .B(n1289), .Y(n2602) );
  OAI21X1 U573 ( .A(n1321), .B(n1288), .C(n2603), .Y(n3747) );
  NAND2X1 U574 ( .A(arr[270]), .B(n1289), .Y(n2603) );
  OAI21X1 U575 ( .A(n1320), .B(n1288), .C(n2604), .Y(n3748) );
  NAND2X1 U576 ( .A(arr[271]), .B(n1289), .Y(n2604) );
  OAI21X1 U578 ( .A(n1335), .B(n1286), .C(n2607), .Y(n3749) );
  NAND2X1 U579 ( .A(arr[272]), .B(n1287), .Y(n2607) );
  OAI21X1 U580 ( .A(n1334), .B(n1286), .C(n2608), .Y(n3750) );
  NAND2X1 U581 ( .A(arr[273]), .B(n1287), .Y(n2608) );
  OAI21X1 U582 ( .A(n1333), .B(n1286), .C(n2609), .Y(n3751) );
  NAND2X1 U583 ( .A(arr[274]), .B(n1286), .Y(n2609) );
  OAI21X1 U584 ( .A(n1332), .B(n1286), .C(n2610), .Y(n3752) );
  NAND2X1 U585 ( .A(arr[275]), .B(n1286), .Y(n2610) );
  OAI21X1 U586 ( .A(n1331), .B(n1286), .C(n2611), .Y(n3753) );
  NAND2X1 U587 ( .A(arr[276]), .B(n1287), .Y(n2611) );
  OAI21X1 U588 ( .A(n1330), .B(n1286), .C(n2612), .Y(n3754) );
  NAND2X1 U589 ( .A(arr[277]), .B(n1287), .Y(n2612) );
  OAI21X1 U590 ( .A(n1329), .B(n1286), .C(n2613), .Y(n3755) );
  NAND2X1 U591 ( .A(arr[278]), .B(n1287), .Y(n2613) );
  OAI21X1 U592 ( .A(n1328), .B(n1286), .C(n2614), .Y(n3756) );
  NAND2X1 U593 ( .A(arr[279]), .B(n1287), .Y(n2614) );
  OAI21X1 U594 ( .A(n1327), .B(n1286), .C(n2615), .Y(n3757) );
  NAND2X1 U595 ( .A(arr[280]), .B(n1287), .Y(n2615) );
  OAI21X1 U596 ( .A(n2309), .B(n1287), .C(n2616), .Y(n3758) );
  NAND2X1 U597 ( .A(arr[281]), .B(n1287), .Y(n2616) );
  OAI21X1 U598 ( .A(n2311), .B(n1287), .C(n2617), .Y(n3759) );
  NAND2X1 U599 ( .A(arr[282]), .B(n1287), .Y(n2617) );
  OAI21X1 U600 ( .A(n2313), .B(n1287), .C(n2618), .Y(n3760) );
  NAND2X1 U601 ( .A(arr[283]), .B(n1287), .Y(n2618) );
  OAI21X1 U602 ( .A(n1323), .B(n1286), .C(n2619), .Y(n3761) );
  NAND2X1 U603 ( .A(arr[284]), .B(n1287), .Y(n2619) );
  OAI21X1 U604 ( .A(n1322), .B(n1286), .C(n2620), .Y(n3762) );
  NAND2X1 U605 ( .A(arr[285]), .B(n1287), .Y(n2620) );
  OAI21X1 U606 ( .A(n1321), .B(n1286), .C(n2621), .Y(n3763) );
  NAND2X1 U607 ( .A(arr[286]), .B(n1287), .Y(n2621) );
  OAI21X1 U608 ( .A(n1320), .B(n1286), .C(n2622), .Y(n3764) );
  NAND2X1 U609 ( .A(arr[287]), .B(n1287), .Y(n2622) );
  OAI21X1 U611 ( .A(n1335), .B(n1284), .C(n2624), .Y(n3765) );
  NAND2X1 U612 ( .A(arr[288]), .B(n1285), .Y(n2624) );
  OAI21X1 U613 ( .A(n1334), .B(n1284), .C(n2625), .Y(n3766) );
  NAND2X1 U614 ( .A(arr[289]), .B(n1285), .Y(n2625) );
  OAI21X1 U615 ( .A(n1333), .B(n1284), .C(n2626), .Y(n3767) );
  NAND2X1 U616 ( .A(arr[290]), .B(n1284), .Y(n2626) );
  OAI21X1 U617 ( .A(n1332), .B(n1284), .C(n2627), .Y(n3768) );
  NAND2X1 U618 ( .A(arr[291]), .B(n1284), .Y(n2627) );
  OAI21X1 U619 ( .A(n1331), .B(n1284), .C(n2628), .Y(n3769) );
  NAND2X1 U620 ( .A(arr[292]), .B(n1285), .Y(n2628) );
  OAI21X1 U621 ( .A(n1330), .B(n1284), .C(n2629), .Y(n3770) );
  NAND2X1 U622 ( .A(arr[293]), .B(n1285), .Y(n2629) );
  OAI21X1 U623 ( .A(n1329), .B(n1284), .C(n2630), .Y(n3771) );
  NAND2X1 U624 ( .A(arr[294]), .B(n1285), .Y(n2630) );
  OAI21X1 U625 ( .A(n1328), .B(n1284), .C(n2631), .Y(n3772) );
  NAND2X1 U626 ( .A(arr[295]), .B(n1285), .Y(n2631) );
  OAI21X1 U627 ( .A(n1327), .B(n1284), .C(n2632), .Y(n3773) );
  NAND2X1 U628 ( .A(arr[296]), .B(n1285), .Y(n2632) );
  OAI21X1 U629 ( .A(n1326), .B(n1285), .C(n2633), .Y(n3774) );
  NAND2X1 U630 ( .A(arr[297]), .B(n1285), .Y(n2633) );
  OAI21X1 U631 ( .A(n1325), .B(n1285), .C(n2634), .Y(n3775) );
  NAND2X1 U632 ( .A(arr[298]), .B(n1285), .Y(n2634) );
  OAI21X1 U633 ( .A(n1324), .B(n1285), .C(n2635), .Y(n3776) );
  NAND2X1 U634 ( .A(arr[299]), .B(n1285), .Y(n2635) );
  OAI21X1 U635 ( .A(n1323), .B(n1284), .C(n2636), .Y(n3777) );
  NAND2X1 U636 ( .A(arr[300]), .B(n1285), .Y(n2636) );
  OAI21X1 U637 ( .A(n1322), .B(n1284), .C(n2637), .Y(n3778) );
  NAND2X1 U638 ( .A(arr[301]), .B(n1285), .Y(n2637) );
  OAI21X1 U639 ( .A(n1321), .B(n1284), .C(n2638), .Y(n3779) );
  NAND2X1 U640 ( .A(arr[302]), .B(n1285), .Y(n2638) );
  OAI21X1 U641 ( .A(n1320), .B(n1284), .C(n2639), .Y(n3780) );
  NAND2X1 U642 ( .A(arr[303]), .B(n1285), .Y(n2639) );
  OAI21X1 U644 ( .A(n1335), .B(n1282), .C(n2642), .Y(n3781) );
  NAND2X1 U645 ( .A(arr[304]), .B(n1283), .Y(n2642) );
  OAI21X1 U646 ( .A(n1334), .B(n1282), .C(n2643), .Y(n3782) );
  NAND2X1 U647 ( .A(arr[305]), .B(n1283), .Y(n2643) );
  OAI21X1 U648 ( .A(n1333), .B(n1282), .C(n2644), .Y(n3783) );
  NAND2X1 U649 ( .A(arr[306]), .B(n1282), .Y(n2644) );
  OAI21X1 U650 ( .A(n1332), .B(n1282), .C(n2645), .Y(n3784) );
  NAND2X1 U651 ( .A(arr[307]), .B(n1282), .Y(n2645) );
  OAI21X1 U652 ( .A(n1331), .B(n1282), .C(n2646), .Y(n3785) );
  NAND2X1 U653 ( .A(arr[308]), .B(n1283), .Y(n2646) );
  OAI21X1 U654 ( .A(n1330), .B(n1282), .C(n2647), .Y(n3786) );
  NAND2X1 U655 ( .A(arr[309]), .B(n1283), .Y(n2647) );
  OAI21X1 U656 ( .A(n1329), .B(n1282), .C(n2648), .Y(n3787) );
  NAND2X1 U657 ( .A(arr[310]), .B(n1283), .Y(n2648) );
  OAI21X1 U658 ( .A(n1328), .B(n1282), .C(n2649), .Y(n3788) );
  NAND2X1 U659 ( .A(arr[311]), .B(n1283), .Y(n2649) );
  OAI21X1 U660 ( .A(n1327), .B(n1282), .C(n2650), .Y(n3789) );
  NAND2X1 U661 ( .A(arr[312]), .B(n1283), .Y(n2650) );
  OAI21X1 U662 ( .A(n1326), .B(n1283), .C(n2651), .Y(n3790) );
  NAND2X1 U663 ( .A(arr[313]), .B(n1283), .Y(n2651) );
  OAI21X1 U664 ( .A(n1325), .B(n1283), .C(n2652), .Y(n3791) );
  NAND2X1 U665 ( .A(arr[314]), .B(n1283), .Y(n2652) );
  OAI21X1 U666 ( .A(n1324), .B(n1283), .C(n2653), .Y(n3792) );
  NAND2X1 U667 ( .A(arr[315]), .B(n1283), .Y(n2653) );
  OAI21X1 U668 ( .A(n1323), .B(n1282), .C(n2654), .Y(n3793) );
  NAND2X1 U669 ( .A(arr[316]), .B(n1283), .Y(n2654) );
  OAI21X1 U670 ( .A(n1322), .B(n1282), .C(n2655), .Y(n3794) );
  NAND2X1 U671 ( .A(arr[317]), .B(n1283), .Y(n2655) );
  OAI21X1 U672 ( .A(n1321), .B(n1282), .C(n2656), .Y(n3795) );
  NAND2X1 U673 ( .A(arr[318]), .B(n1283), .Y(n2656) );
  OAI21X1 U674 ( .A(n1320), .B(n1282), .C(n2657), .Y(n3796) );
  NAND2X1 U675 ( .A(arr[319]), .B(n1283), .Y(n2657) );
  OAI21X1 U677 ( .A(n1335), .B(n1280), .C(n2659), .Y(n3797) );
  NAND2X1 U678 ( .A(arr[320]), .B(n1281), .Y(n2659) );
  OAI21X1 U679 ( .A(n1334), .B(n1280), .C(n2660), .Y(n3798) );
  NAND2X1 U680 ( .A(arr[321]), .B(n1281), .Y(n2660) );
  OAI21X1 U681 ( .A(n1333), .B(n1280), .C(n2661), .Y(n3799) );
  NAND2X1 U682 ( .A(arr[322]), .B(n1280), .Y(n2661) );
  OAI21X1 U683 ( .A(n1332), .B(n1280), .C(n2662), .Y(n3800) );
  NAND2X1 U684 ( .A(arr[323]), .B(n1280), .Y(n2662) );
  OAI21X1 U685 ( .A(n1331), .B(n1280), .C(n2663), .Y(n3801) );
  NAND2X1 U686 ( .A(arr[324]), .B(n1281), .Y(n2663) );
  OAI21X1 U687 ( .A(n1330), .B(n1280), .C(n2664), .Y(n3802) );
  NAND2X1 U688 ( .A(arr[325]), .B(n1281), .Y(n2664) );
  OAI21X1 U689 ( .A(n1329), .B(n1280), .C(n2665), .Y(n3803) );
  NAND2X1 U690 ( .A(arr[326]), .B(n1281), .Y(n2665) );
  OAI21X1 U691 ( .A(n1328), .B(n1280), .C(n2666), .Y(n3804) );
  NAND2X1 U692 ( .A(arr[327]), .B(n1281), .Y(n2666) );
  OAI21X1 U693 ( .A(n1327), .B(n1280), .C(n2667), .Y(n3805) );
  NAND2X1 U694 ( .A(arr[328]), .B(n1281), .Y(n2667) );
  OAI21X1 U695 ( .A(n1326), .B(n1281), .C(n2668), .Y(n3806) );
  NAND2X1 U696 ( .A(arr[329]), .B(n1281), .Y(n2668) );
  OAI21X1 U697 ( .A(n1325), .B(n1281), .C(n2669), .Y(n3807) );
  NAND2X1 U698 ( .A(arr[330]), .B(n1281), .Y(n2669) );
  OAI21X1 U699 ( .A(n1324), .B(n1281), .C(n2670), .Y(n3808) );
  NAND2X1 U700 ( .A(arr[331]), .B(n1281), .Y(n2670) );
  OAI21X1 U701 ( .A(n1323), .B(n1280), .C(n2671), .Y(n3809) );
  NAND2X1 U702 ( .A(arr[332]), .B(n1281), .Y(n2671) );
  OAI21X1 U703 ( .A(n1322), .B(n1280), .C(n2672), .Y(n3810) );
  NAND2X1 U704 ( .A(arr[333]), .B(n1281), .Y(n2672) );
  OAI21X1 U705 ( .A(n1321), .B(n1280), .C(n2673), .Y(n3811) );
  NAND2X1 U706 ( .A(arr[334]), .B(n1281), .Y(n2673) );
  OAI21X1 U707 ( .A(n1320), .B(n1280), .C(n2674), .Y(n3812) );
  NAND2X1 U708 ( .A(arr[335]), .B(n1281), .Y(n2674) );
  OAI21X1 U710 ( .A(n1335), .B(n1278), .C(n2677), .Y(n3813) );
  NAND2X1 U711 ( .A(arr[336]), .B(n1279), .Y(n2677) );
  OAI21X1 U712 ( .A(n1334), .B(n1278), .C(n2678), .Y(n3814) );
  NAND2X1 U713 ( .A(arr[337]), .B(n1279), .Y(n2678) );
  OAI21X1 U714 ( .A(n1333), .B(n1278), .C(n2679), .Y(n3815) );
  NAND2X1 U715 ( .A(arr[338]), .B(n1278), .Y(n2679) );
  OAI21X1 U716 ( .A(n1332), .B(n1278), .C(n2680), .Y(n3816) );
  NAND2X1 U717 ( .A(arr[339]), .B(n1278), .Y(n2680) );
  OAI21X1 U718 ( .A(n1331), .B(n1278), .C(n2681), .Y(n3817) );
  NAND2X1 U719 ( .A(arr[340]), .B(n1279), .Y(n2681) );
  OAI21X1 U720 ( .A(n1330), .B(n1278), .C(n2682), .Y(n3818) );
  NAND2X1 U721 ( .A(arr[341]), .B(n1279), .Y(n2682) );
  OAI21X1 U722 ( .A(n1329), .B(n1278), .C(n2683), .Y(n3819) );
  NAND2X1 U723 ( .A(arr[342]), .B(n1279), .Y(n2683) );
  OAI21X1 U724 ( .A(n1328), .B(n1278), .C(n2684), .Y(n3820) );
  NAND2X1 U725 ( .A(arr[343]), .B(n1279), .Y(n2684) );
  OAI21X1 U726 ( .A(n1327), .B(n1278), .C(n2685), .Y(n3821) );
  NAND2X1 U727 ( .A(arr[344]), .B(n1279), .Y(n2685) );
  OAI21X1 U728 ( .A(n1326), .B(n1279), .C(n2686), .Y(n3822) );
  NAND2X1 U729 ( .A(arr[345]), .B(n1279), .Y(n2686) );
  OAI21X1 U730 ( .A(n1325), .B(n1279), .C(n2687), .Y(n3823) );
  NAND2X1 U731 ( .A(arr[346]), .B(n1279), .Y(n2687) );
  OAI21X1 U732 ( .A(n1324), .B(n1279), .C(n2688), .Y(n3824) );
  NAND2X1 U733 ( .A(arr[347]), .B(n1279), .Y(n2688) );
  OAI21X1 U734 ( .A(n1323), .B(n1278), .C(n2689), .Y(n3825) );
  NAND2X1 U735 ( .A(arr[348]), .B(n1279), .Y(n2689) );
  OAI21X1 U736 ( .A(n1322), .B(n1278), .C(n2690), .Y(n3826) );
  NAND2X1 U737 ( .A(arr[349]), .B(n1279), .Y(n2690) );
  OAI21X1 U738 ( .A(n1321), .B(n1278), .C(n2691), .Y(n3827) );
  NAND2X1 U739 ( .A(arr[350]), .B(n1279), .Y(n2691) );
  OAI21X1 U740 ( .A(n1320), .B(n1278), .C(n2692), .Y(n3828) );
  NAND2X1 U741 ( .A(arr[351]), .B(n1279), .Y(n2692) );
  OAI21X1 U743 ( .A(n1335), .B(n1276), .C(n2694), .Y(n3829) );
  NAND2X1 U744 ( .A(arr[352]), .B(n1277), .Y(n2694) );
  OAI21X1 U745 ( .A(n1334), .B(n1276), .C(n2695), .Y(n3830) );
  NAND2X1 U746 ( .A(arr[353]), .B(n1277), .Y(n2695) );
  OAI21X1 U747 ( .A(n1333), .B(n1276), .C(n2696), .Y(n3831) );
  NAND2X1 U748 ( .A(arr[354]), .B(n1276), .Y(n2696) );
  OAI21X1 U749 ( .A(n1332), .B(n1276), .C(n2697), .Y(n3832) );
  NAND2X1 U750 ( .A(arr[355]), .B(n1276), .Y(n2697) );
  OAI21X1 U751 ( .A(n1331), .B(n1276), .C(n2698), .Y(n3833) );
  NAND2X1 U752 ( .A(arr[356]), .B(n1277), .Y(n2698) );
  OAI21X1 U753 ( .A(n1330), .B(n1276), .C(n2699), .Y(n3834) );
  NAND2X1 U754 ( .A(arr[357]), .B(n1277), .Y(n2699) );
  OAI21X1 U755 ( .A(n1329), .B(n1276), .C(n2700), .Y(n3835) );
  NAND2X1 U756 ( .A(arr[358]), .B(n1277), .Y(n2700) );
  OAI21X1 U757 ( .A(n1328), .B(n1276), .C(n2701), .Y(n3836) );
  NAND2X1 U758 ( .A(arr[359]), .B(n1277), .Y(n2701) );
  OAI21X1 U759 ( .A(n1327), .B(n1276), .C(n2702), .Y(n3837) );
  NAND2X1 U760 ( .A(arr[360]), .B(n1277), .Y(n2702) );
  OAI21X1 U761 ( .A(n1326), .B(n1277), .C(n2703), .Y(n3838) );
  NAND2X1 U762 ( .A(arr[361]), .B(n1277), .Y(n2703) );
  OAI21X1 U763 ( .A(n1325), .B(n1277), .C(n2704), .Y(n3839) );
  NAND2X1 U764 ( .A(arr[362]), .B(n1277), .Y(n2704) );
  OAI21X1 U765 ( .A(n1324), .B(n1277), .C(n2705), .Y(n3840) );
  NAND2X1 U766 ( .A(arr[363]), .B(n1277), .Y(n2705) );
  OAI21X1 U767 ( .A(n1323), .B(n1276), .C(n2706), .Y(n3841) );
  NAND2X1 U768 ( .A(arr[364]), .B(n1277), .Y(n2706) );
  OAI21X1 U769 ( .A(n1322), .B(n1276), .C(n2707), .Y(n3842) );
  NAND2X1 U770 ( .A(arr[365]), .B(n1277), .Y(n2707) );
  OAI21X1 U771 ( .A(n1321), .B(n1276), .C(n2708), .Y(n3843) );
  NAND2X1 U772 ( .A(arr[366]), .B(n1277), .Y(n2708) );
  OAI21X1 U773 ( .A(n1320), .B(n1276), .C(n2709), .Y(n3844) );
  NAND2X1 U774 ( .A(arr[367]), .B(n1277), .Y(n2709) );
  OAI21X1 U776 ( .A(n2291), .B(n1274), .C(n2712), .Y(n3845) );
  NAND2X1 U777 ( .A(arr[368]), .B(n1275), .Y(n2712) );
  OAI21X1 U778 ( .A(n2293), .B(n1274), .C(n2713), .Y(n3846) );
  NAND2X1 U779 ( .A(arr[369]), .B(n1275), .Y(n2713) );
  OAI21X1 U780 ( .A(n2295), .B(n1274), .C(n2714), .Y(n3847) );
  NAND2X1 U781 ( .A(arr[370]), .B(n1274), .Y(n2714) );
  OAI21X1 U782 ( .A(n2297), .B(n1274), .C(n2715), .Y(n3848) );
  NAND2X1 U783 ( .A(arr[371]), .B(n1274), .Y(n2715) );
  OAI21X1 U784 ( .A(n2299), .B(n1274), .C(n2716), .Y(n3849) );
  NAND2X1 U785 ( .A(arr[372]), .B(n1275), .Y(n2716) );
  OAI21X1 U786 ( .A(n2301), .B(n1274), .C(n2717), .Y(n3850) );
  NAND2X1 U787 ( .A(arr[373]), .B(n1275), .Y(n2717) );
  OAI21X1 U788 ( .A(n2303), .B(n1274), .C(n2718), .Y(n3851) );
  NAND2X1 U789 ( .A(arr[374]), .B(n1275), .Y(n2718) );
  OAI21X1 U790 ( .A(n2305), .B(n1274), .C(n2719), .Y(n3852) );
  NAND2X1 U791 ( .A(arr[375]), .B(n1275), .Y(n2719) );
  OAI21X1 U792 ( .A(n2307), .B(n1274), .C(n2720), .Y(n3853) );
  NAND2X1 U793 ( .A(arr[376]), .B(n1275), .Y(n2720) );
  OAI21X1 U794 ( .A(n2309), .B(n1275), .C(n2721), .Y(n3854) );
  NAND2X1 U795 ( .A(arr[377]), .B(n1275), .Y(n2721) );
  OAI21X1 U796 ( .A(n2311), .B(n1275), .C(n2722), .Y(n3855) );
  NAND2X1 U797 ( .A(arr[378]), .B(n1275), .Y(n2722) );
  OAI21X1 U798 ( .A(n2313), .B(n1275), .C(n2723), .Y(n3856) );
  NAND2X1 U799 ( .A(arr[379]), .B(n1275), .Y(n2723) );
  OAI21X1 U800 ( .A(n2315), .B(n1274), .C(n2724), .Y(n3857) );
  NAND2X1 U801 ( .A(arr[380]), .B(n1275), .Y(n2724) );
  OAI21X1 U802 ( .A(n2317), .B(n1274), .C(n2725), .Y(n3858) );
  NAND2X1 U803 ( .A(arr[381]), .B(n1275), .Y(n2725) );
  OAI21X1 U804 ( .A(n2319), .B(n1274), .C(n2726), .Y(n3859) );
  NAND2X1 U805 ( .A(arr[382]), .B(n1275), .Y(n2726) );
  OAI21X1 U806 ( .A(n2321), .B(n1274), .C(n2727), .Y(n3860) );
  NAND2X1 U807 ( .A(arr[383]), .B(n1275), .Y(n2727) );
  OAI21X1 U809 ( .A(n1335), .B(n1272), .C(n2729), .Y(n3861) );
  NAND2X1 U810 ( .A(arr[384]), .B(n1273), .Y(n2729) );
  OAI21X1 U811 ( .A(n1334), .B(n1272), .C(n2730), .Y(n3862) );
  NAND2X1 U812 ( .A(arr[385]), .B(n1273), .Y(n2730) );
  OAI21X1 U813 ( .A(n1333), .B(n1272), .C(n2731), .Y(n3863) );
  NAND2X1 U814 ( .A(arr[386]), .B(n1272), .Y(n2731) );
  OAI21X1 U815 ( .A(n1332), .B(n1272), .C(n2732), .Y(n3864) );
  NAND2X1 U816 ( .A(arr[387]), .B(n1272), .Y(n2732) );
  OAI21X1 U817 ( .A(n1331), .B(n1272), .C(n2733), .Y(n3865) );
  NAND2X1 U818 ( .A(arr[388]), .B(n1273), .Y(n2733) );
  OAI21X1 U819 ( .A(n1330), .B(n1272), .C(n2734), .Y(n3866) );
  NAND2X1 U820 ( .A(arr[389]), .B(n1273), .Y(n2734) );
  OAI21X1 U821 ( .A(n1329), .B(n1272), .C(n2735), .Y(n3867) );
  NAND2X1 U822 ( .A(arr[390]), .B(n1273), .Y(n2735) );
  OAI21X1 U823 ( .A(n1328), .B(n1272), .C(n2736), .Y(n3868) );
  NAND2X1 U824 ( .A(arr[391]), .B(n1273), .Y(n2736) );
  OAI21X1 U825 ( .A(n1327), .B(n1272), .C(n2737), .Y(n3869) );
  NAND2X1 U826 ( .A(arr[392]), .B(n1273), .Y(n2737) );
  OAI21X1 U827 ( .A(n1326), .B(n1273), .C(n2738), .Y(n3870) );
  NAND2X1 U828 ( .A(arr[393]), .B(n1273), .Y(n2738) );
  OAI21X1 U829 ( .A(n1325), .B(n1273), .C(n2739), .Y(n3871) );
  NAND2X1 U830 ( .A(arr[394]), .B(n1273), .Y(n2739) );
  OAI21X1 U831 ( .A(n1324), .B(n1273), .C(n2740), .Y(n3872) );
  NAND2X1 U832 ( .A(arr[395]), .B(n1273), .Y(n2740) );
  OAI21X1 U833 ( .A(n1323), .B(n1272), .C(n2741), .Y(n3873) );
  NAND2X1 U834 ( .A(arr[396]), .B(n1273), .Y(n2741) );
  OAI21X1 U835 ( .A(n1322), .B(n1272), .C(n2742), .Y(n3874) );
  NAND2X1 U836 ( .A(arr[397]), .B(n1273), .Y(n2742) );
  OAI21X1 U837 ( .A(n1321), .B(n1272), .C(n2743), .Y(n3875) );
  NAND2X1 U838 ( .A(arr[398]), .B(n1273), .Y(n2743) );
  OAI21X1 U839 ( .A(n1320), .B(n1272), .C(n2744), .Y(n3876) );
  NAND2X1 U840 ( .A(arr[399]), .B(n1273), .Y(n2744) );
  OAI21X1 U842 ( .A(n2291), .B(n1270), .C(n2747), .Y(n3877) );
  NAND2X1 U843 ( .A(arr[400]), .B(n1271), .Y(n2747) );
  OAI21X1 U844 ( .A(n2293), .B(n1270), .C(n2748), .Y(n3878) );
  NAND2X1 U845 ( .A(arr[401]), .B(n1271), .Y(n2748) );
  OAI21X1 U846 ( .A(n2295), .B(n1270), .C(n2749), .Y(n3879) );
  NAND2X1 U847 ( .A(arr[402]), .B(n1270), .Y(n2749) );
  OAI21X1 U848 ( .A(n2297), .B(n1270), .C(n2750), .Y(n3880) );
  NAND2X1 U849 ( .A(arr[403]), .B(n1270), .Y(n2750) );
  OAI21X1 U850 ( .A(n2299), .B(n1270), .C(n2751), .Y(n3881) );
  NAND2X1 U851 ( .A(arr[404]), .B(n1271), .Y(n2751) );
  OAI21X1 U852 ( .A(n2301), .B(n1270), .C(n2752), .Y(n3882) );
  NAND2X1 U853 ( .A(arr[405]), .B(n1271), .Y(n2752) );
  OAI21X1 U854 ( .A(n2303), .B(n1270), .C(n2753), .Y(n3883) );
  NAND2X1 U855 ( .A(arr[406]), .B(n1271), .Y(n2753) );
  OAI21X1 U856 ( .A(n2305), .B(n1270), .C(n2754), .Y(n3884) );
  NAND2X1 U857 ( .A(arr[407]), .B(n1271), .Y(n2754) );
  OAI21X1 U858 ( .A(n2307), .B(n1270), .C(n2755), .Y(n3885) );
  NAND2X1 U859 ( .A(arr[408]), .B(n1271), .Y(n2755) );
  OAI21X1 U860 ( .A(n1326), .B(n1271), .C(n2756), .Y(n3886) );
  NAND2X1 U861 ( .A(arr[409]), .B(n1271), .Y(n2756) );
  OAI21X1 U862 ( .A(n1325), .B(n1271), .C(n2757), .Y(n3887) );
  NAND2X1 U863 ( .A(arr[410]), .B(n1271), .Y(n2757) );
  OAI21X1 U864 ( .A(n1324), .B(n1271), .C(n2758), .Y(n3888) );
  NAND2X1 U865 ( .A(arr[411]), .B(n1271), .Y(n2758) );
  OAI21X1 U866 ( .A(n2315), .B(n1270), .C(n2759), .Y(n3889) );
  NAND2X1 U867 ( .A(arr[412]), .B(n1271), .Y(n2759) );
  OAI21X1 U868 ( .A(n2317), .B(n1270), .C(n2760), .Y(n3890) );
  NAND2X1 U869 ( .A(arr[413]), .B(n1271), .Y(n2760) );
  OAI21X1 U870 ( .A(n2319), .B(n1270), .C(n2761), .Y(n3891) );
  NAND2X1 U871 ( .A(arr[414]), .B(n1271), .Y(n2761) );
  OAI21X1 U872 ( .A(n2321), .B(n1270), .C(n2762), .Y(n3892) );
  NAND2X1 U873 ( .A(arr[415]), .B(n1271), .Y(n2762) );
  OAI21X1 U875 ( .A(n2291), .B(n1268), .C(n2764), .Y(n3893) );
  NAND2X1 U876 ( .A(arr[416]), .B(n1269), .Y(n2764) );
  OAI21X1 U877 ( .A(n2293), .B(n1268), .C(n2765), .Y(n3894) );
  NAND2X1 U878 ( .A(arr[417]), .B(n1269), .Y(n2765) );
  OAI21X1 U879 ( .A(n2295), .B(n1268), .C(n2766), .Y(n3895) );
  NAND2X1 U880 ( .A(arr[418]), .B(n1268), .Y(n2766) );
  OAI21X1 U881 ( .A(n2297), .B(n1268), .C(n2767), .Y(n3896) );
  NAND2X1 U882 ( .A(arr[419]), .B(n1268), .Y(n2767) );
  OAI21X1 U883 ( .A(n2299), .B(n1268), .C(n2768), .Y(n3897) );
  NAND2X1 U884 ( .A(arr[420]), .B(n1269), .Y(n2768) );
  OAI21X1 U885 ( .A(n2301), .B(n1268), .C(n2769), .Y(n3898) );
  NAND2X1 U886 ( .A(arr[421]), .B(n1269), .Y(n2769) );
  OAI21X1 U887 ( .A(n2303), .B(n1268), .C(n2770), .Y(n3899) );
  NAND2X1 U888 ( .A(arr[422]), .B(n1269), .Y(n2770) );
  OAI21X1 U889 ( .A(n2305), .B(n1268), .C(n2771), .Y(n3900) );
  NAND2X1 U890 ( .A(arr[423]), .B(n1269), .Y(n2771) );
  OAI21X1 U891 ( .A(n2307), .B(n1268), .C(n2772), .Y(n3901) );
  NAND2X1 U892 ( .A(arr[424]), .B(n1269), .Y(n2772) );
  OAI21X1 U893 ( .A(n2309), .B(n1269), .C(n2773), .Y(n3902) );
  NAND2X1 U894 ( .A(arr[425]), .B(n1269), .Y(n2773) );
  OAI21X1 U895 ( .A(n2311), .B(n1269), .C(n2774), .Y(n3903) );
  NAND2X1 U896 ( .A(arr[426]), .B(n1269), .Y(n2774) );
  OAI21X1 U897 ( .A(n2313), .B(n1269), .C(n2775), .Y(n3904) );
  NAND2X1 U898 ( .A(arr[427]), .B(n1269), .Y(n2775) );
  OAI21X1 U899 ( .A(n2315), .B(n1268), .C(n2776), .Y(n3905) );
  NAND2X1 U900 ( .A(arr[428]), .B(n1269), .Y(n2776) );
  OAI21X1 U901 ( .A(n2317), .B(n1268), .C(n2777), .Y(n3906) );
  NAND2X1 U902 ( .A(arr[429]), .B(n1269), .Y(n2777) );
  OAI21X1 U903 ( .A(n2319), .B(n1268), .C(n2778), .Y(n3907) );
  NAND2X1 U904 ( .A(arr[430]), .B(n1269), .Y(n2778) );
  OAI21X1 U905 ( .A(n2321), .B(n1268), .C(n2779), .Y(n3908) );
  NAND2X1 U906 ( .A(arr[431]), .B(n1269), .Y(n2779) );
  OAI21X1 U908 ( .A(n2291), .B(n1266), .C(n2782), .Y(n3909) );
  NAND2X1 U909 ( .A(arr[432]), .B(n1267), .Y(n2782) );
  OAI21X1 U910 ( .A(n2293), .B(n1266), .C(n2783), .Y(n3910) );
  NAND2X1 U911 ( .A(arr[433]), .B(n1267), .Y(n2783) );
  OAI21X1 U912 ( .A(n2295), .B(n1266), .C(n2784), .Y(n3911) );
  NAND2X1 U913 ( .A(arr[434]), .B(n1266), .Y(n2784) );
  OAI21X1 U914 ( .A(n2297), .B(n1266), .C(n2785), .Y(n3912) );
  NAND2X1 U915 ( .A(arr[435]), .B(n1266), .Y(n2785) );
  OAI21X1 U916 ( .A(n2299), .B(n1266), .C(n2786), .Y(n3913) );
  NAND2X1 U917 ( .A(arr[436]), .B(n1267), .Y(n2786) );
  OAI21X1 U918 ( .A(n2301), .B(n1266), .C(n2787), .Y(n3914) );
  NAND2X1 U919 ( .A(arr[437]), .B(n1267), .Y(n2787) );
  OAI21X1 U920 ( .A(n2303), .B(n1266), .C(n2788), .Y(n3915) );
  NAND2X1 U921 ( .A(arr[438]), .B(n1267), .Y(n2788) );
  OAI21X1 U922 ( .A(n2305), .B(n1266), .C(n2789), .Y(n3916) );
  NAND2X1 U923 ( .A(arr[439]), .B(n1267), .Y(n2789) );
  OAI21X1 U924 ( .A(n2307), .B(n1266), .C(n2790), .Y(n3917) );
  NAND2X1 U925 ( .A(arr[440]), .B(n1267), .Y(n2790) );
  OAI21X1 U926 ( .A(n2309), .B(n1267), .C(n2791), .Y(n3918) );
  NAND2X1 U927 ( .A(arr[441]), .B(n1267), .Y(n2791) );
  OAI21X1 U928 ( .A(n2311), .B(n1267), .C(n2792), .Y(n3919) );
  NAND2X1 U929 ( .A(arr[442]), .B(n1267), .Y(n2792) );
  OAI21X1 U930 ( .A(n2313), .B(n1267), .C(n2793), .Y(n3920) );
  NAND2X1 U931 ( .A(arr[443]), .B(n1267), .Y(n2793) );
  OAI21X1 U932 ( .A(n2315), .B(n1266), .C(n2794), .Y(n3921) );
  NAND2X1 U933 ( .A(arr[444]), .B(n1267), .Y(n2794) );
  OAI21X1 U934 ( .A(n2317), .B(n1266), .C(n2795), .Y(n3922) );
  NAND2X1 U935 ( .A(arr[445]), .B(n1267), .Y(n2795) );
  OAI21X1 U936 ( .A(n2319), .B(n1266), .C(n2796), .Y(n3923) );
  NAND2X1 U937 ( .A(arr[446]), .B(n1267), .Y(n2796) );
  OAI21X1 U938 ( .A(n2321), .B(n1266), .C(n2797), .Y(n3924) );
  NAND2X1 U939 ( .A(arr[447]), .B(n1267), .Y(n2797) );
  OAI21X1 U941 ( .A(n2291), .B(n1264), .C(n2799), .Y(n3925) );
  NAND2X1 U942 ( .A(arr[448]), .B(n1265), .Y(n2799) );
  OAI21X1 U943 ( .A(n2293), .B(n1264), .C(n2800), .Y(n3926) );
  NAND2X1 U944 ( .A(arr[449]), .B(n1265), .Y(n2800) );
  OAI21X1 U945 ( .A(n2295), .B(n1264), .C(n2801), .Y(n3927) );
  NAND2X1 U946 ( .A(arr[450]), .B(n1264), .Y(n2801) );
  OAI21X1 U947 ( .A(n2297), .B(n1264), .C(n2802), .Y(n3928) );
  NAND2X1 U948 ( .A(arr[451]), .B(n1264), .Y(n2802) );
  OAI21X1 U949 ( .A(n2299), .B(n1264), .C(n2803), .Y(n3929) );
  NAND2X1 U950 ( .A(arr[452]), .B(n1265), .Y(n2803) );
  OAI21X1 U951 ( .A(n2301), .B(n1264), .C(n2804), .Y(n3930) );
  NAND2X1 U952 ( .A(arr[453]), .B(n1265), .Y(n2804) );
  OAI21X1 U953 ( .A(n2303), .B(n1264), .C(n2805), .Y(n3931) );
  NAND2X1 U954 ( .A(arr[454]), .B(n1265), .Y(n2805) );
  OAI21X1 U955 ( .A(n2305), .B(n1264), .C(n2806), .Y(n3932) );
  NAND2X1 U956 ( .A(arr[455]), .B(n1265), .Y(n2806) );
  OAI21X1 U957 ( .A(n2307), .B(n1264), .C(n2807), .Y(n3933) );
  NAND2X1 U958 ( .A(arr[456]), .B(n1265), .Y(n2807) );
  OAI21X1 U959 ( .A(n2309), .B(n1265), .C(n2808), .Y(n3934) );
  NAND2X1 U960 ( .A(arr[457]), .B(n1265), .Y(n2808) );
  OAI21X1 U961 ( .A(n2311), .B(n1265), .C(n2809), .Y(n3935) );
  NAND2X1 U962 ( .A(arr[458]), .B(n1265), .Y(n2809) );
  OAI21X1 U963 ( .A(n2313), .B(n1265), .C(n2810), .Y(n3936) );
  NAND2X1 U964 ( .A(arr[459]), .B(n1265), .Y(n2810) );
  OAI21X1 U965 ( .A(n2315), .B(n1264), .C(n2811), .Y(n3937) );
  NAND2X1 U966 ( .A(arr[460]), .B(n1265), .Y(n2811) );
  OAI21X1 U967 ( .A(n2317), .B(n1264), .C(n2812), .Y(n3938) );
  NAND2X1 U968 ( .A(arr[461]), .B(n1265), .Y(n2812) );
  OAI21X1 U969 ( .A(n2319), .B(n1264), .C(n2813), .Y(n3939) );
  NAND2X1 U970 ( .A(arr[462]), .B(n1265), .Y(n2813) );
  OAI21X1 U971 ( .A(n2321), .B(n1264), .C(n2814), .Y(n3940) );
  NAND2X1 U972 ( .A(arr[463]), .B(n1265), .Y(n2814) );
  OAI21X1 U974 ( .A(n2291), .B(n1262), .C(n2817), .Y(n3941) );
  NAND2X1 U975 ( .A(arr[464]), .B(n1263), .Y(n2817) );
  OAI21X1 U976 ( .A(n2293), .B(n1262), .C(n2818), .Y(n3942) );
  NAND2X1 U977 ( .A(arr[465]), .B(n1263), .Y(n2818) );
  OAI21X1 U978 ( .A(n2295), .B(n1262), .C(n2819), .Y(n3943) );
  NAND2X1 U979 ( .A(arr[466]), .B(n1262), .Y(n2819) );
  OAI21X1 U980 ( .A(n2297), .B(n1262), .C(n2820), .Y(n3944) );
  NAND2X1 U981 ( .A(arr[467]), .B(n1262), .Y(n2820) );
  OAI21X1 U982 ( .A(n2299), .B(n1262), .C(n2821), .Y(n3945) );
  NAND2X1 U983 ( .A(arr[468]), .B(n1263), .Y(n2821) );
  OAI21X1 U984 ( .A(n2301), .B(n1262), .C(n2822), .Y(n3946) );
  NAND2X1 U985 ( .A(arr[469]), .B(n1263), .Y(n2822) );
  OAI21X1 U986 ( .A(n2303), .B(n1262), .C(n2823), .Y(n3947) );
  NAND2X1 U987 ( .A(arr[470]), .B(n1263), .Y(n2823) );
  OAI21X1 U988 ( .A(n2305), .B(n1262), .C(n2824), .Y(n3948) );
  NAND2X1 U989 ( .A(arr[471]), .B(n1263), .Y(n2824) );
  OAI21X1 U990 ( .A(n2307), .B(n1262), .C(n2825), .Y(n3949) );
  NAND2X1 U991 ( .A(arr[472]), .B(n1263), .Y(n2825) );
  OAI21X1 U992 ( .A(n2309), .B(n1263), .C(n2826), .Y(n3950) );
  NAND2X1 U993 ( .A(arr[473]), .B(n1263), .Y(n2826) );
  OAI21X1 U994 ( .A(n2311), .B(n1263), .C(n2827), .Y(n3951) );
  NAND2X1 U995 ( .A(arr[474]), .B(n1263), .Y(n2827) );
  OAI21X1 U996 ( .A(n2313), .B(n1263), .C(n2828), .Y(n3952) );
  NAND2X1 U997 ( .A(arr[475]), .B(n1263), .Y(n2828) );
  OAI21X1 U998 ( .A(n2315), .B(n1262), .C(n2829), .Y(n3953) );
  NAND2X1 U999 ( .A(arr[476]), .B(n1263), .Y(n2829) );
  OAI21X1 U1000 ( .A(n2317), .B(n1262), .C(n2830), .Y(n3954) );
  NAND2X1 U1001 ( .A(arr[477]), .B(n1263), .Y(n2830) );
  OAI21X1 U1002 ( .A(n2319), .B(n1262), .C(n2831), .Y(n3955) );
  NAND2X1 U1003 ( .A(arr[478]), .B(n1263), .Y(n2831) );
  OAI21X1 U1004 ( .A(n2321), .B(n1262), .C(n2832), .Y(n3956) );
  NAND2X1 U1005 ( .A(arr[479]), .B(n1263), .Y(n2832) );
  OAI21X1 U1007 ( .A(n2291), .B(n1260), .C(n2834), .Y(n3957) );
  NAND2X1 U1008 ( .A(arr[480]), .B(n1261), .Y(n2834) );
  OAI21X1 U1009 ( .A(n2293), .B(n1260), .C(n2835), .Y(n3958) );
  NAND2X1 U1010 ( .A(arr[481]), .B(n1261), .Y(n2835) );
  OAI21X1 U1011 ( .A(n2295), .B(n1260), .C(n2836), .Y(n3959) );
  NAND2X1 U1012 ( .A(arr[482]), .B(n1260), .Y(n2836) );
  OAI21X1 U1013 ( .A(n2297), .B(n1260), .C(n2837), .Y(n3960) );
  NAND2X1 U1014 ( .A(arr[483]), .B(n1260), .Y(n2837) );
  OAI21X1 U1015 ( .A(n2299), .B(n1260), .C(n2838), .Y(n3961) );
  NAND2X1 U1016 ( .A(arr[484]), .B(n1261), .Y(n2838) );
  OAI21X1 U1017 ( .A(n2301), .B(n1260), .C(n2839), .Y(n3962) );
  NAND2X1 U1018 ( .A(arr[485]), .B(n1261), .Y(n2839) );
  OAI21X1 U1019 ( .A(n2303), .B(n1260), .C(n2840), .Y(n3963) );
  NAND2X1 U1020 ( .A(arr[486]), .B(n1261), .Y(n2840) );
  OAI21X1 U1021 ( .A(n2305), .B(n1260), .C(n2841), .Y(n3964) );
  NAND2X1 U1022 ( .A(arr[487]), .B(n1261), .Y(n2841) );
  OAI21X1 U1023 ( .A(n2307), .B(n1260), .C(n2842), .Y(n3965) );
  NAND2X1 U1024 ( .A(arr[488]), .B(n1261), .Y(n2842) );
  OAI21X1 U1025 ( .A(n2309), .B(n1261), .C(n2843), .Y(n3966) );
  NAND2X1 U1026 ( .A(arr[489]), .B(n1261), .Y(n2843) );
  OAI21X1 U1027 ( .A(n2311), .B(n1261), .C(n2844), .Y(n3967) );
  NAND2X1 U1028 ( .A(arr[490]), .B(n1261), .Y(n2844) );
  OAI21X1 U1029 ( .A(n2313), .B(n1261), .C(n2845), .Y(n3968) );
  NAND2X1 U1030 ( .A(arr[491]), .B(n1261), .Y(n2845) );
  OAI21X1 U1031 ( .A(n2315), .B(n1260), .C(n2846), .Y(n3969) );
  NAND2X1 U1032 ( .A(arr[492]), .B(n1261), .Y(n2846) );
  OAI21X1 U1033 ( .A(n2317), .B(n1260), .C(n2847), .Y(n3970) );
  NAND2X1 U1034 ( .A(arr[493]), .B(n1261), .Y(n2847) );
  OAI21X1 U1035 ( .A(n2319), .B(n1260), .C(n2848), .Y(n3971) );
  NAND2X1 U1036 ( .A(arr[494]), .B(n1261), .Y(n2848) );
  OAI21X1 U1037 ( .A(n2321), .B(n1260), .C(n2849), .Y(n3972) );
  NAND2X1 U1038 ( .A(arr[495]), .B(n1261), .Y(n2849) );
  OAI21X1 U1041 ( .A(n2291), .B(n1258), .C(n2854), .Y(n3973) );
  NAND2X1 U1042 ( .A(arr[496]), .B(n1259), .Y(n2854) );
  OAI21X1 U1043 ( .A(n2293), .B(n1258), .C(n2855), .Y(n3974) );
  NAND2X1 U1044 ( .A(arr[497]), .B(n1259), .Y(n2855) );
  OAI21X1 U1045 ( .A(n2295), .B(n1258), .C(n2856), .Y(n3975) );
  NAND2X1 U1046 ( .A(arr[498]), .B(n1258), .Y(n2856) );
  OAI21X1 U1047 ( .A(n2297), .B(n1258), .C(n2857), .Y(n3976) );
  NAND2X1 U1048 ( .A(arr[499]), .B(n1258), .Y(n2857) );
  OAI21X1 U1049 ( .A(n2299), .B(n1258), .C(n2858), .Y(n3977) );
  NAND2X1 U1050 ( .A(arr[500]), .B(n1259), .Y(n2858) );
  OAI21X1 U1051 ( .A(n2301), .B(n1258), .C(n2859), .Y(n3978) );
  NAND2X1 U1052 ( .A(arr[501]), .B(n1259), .Y(n2859) );
  OAI21X1 U1053 ( .A(n2303), .B(n1258), .C(n2860), .Y(n3979) );
  NAND2X1 U1054 ( .A(arr[502]), .B(n1259), .Y(n2860) );
  OAI21X1 U1055 ( .A(n2305), .B(n1258), .C(n2861), .Y(n3980) );
  NAND2X1 U1056 ( .A(arr[503]), .B(n1259), .Y(n2861) );
  OAI21X1 U1057 ( .A(n2307), .B(n1258), .C(n2862), .Y(n3981) );
  NAND2X1 U1058 ( .A(arr[504]), .B(n1259), .Y(n2862) );
  OAI21X1 U1059 ( .A(n2309), .B(n1259), .C(n2863), .Y(n3982) );
  NAND2X1 U1060 ( .A(arr[505]), .B(n1259), .Y(n2863) );
  OAI21X1 U1061 ( .A(n2311), .B(n1259), .C(n2864), .Y(n3983) );
  NAND2X1 U1062 ( .A(arr[506]), .B(n1259), .Y(n2864) );
  OAI21X1 U1063 ( .A(n2313), .B(n1259), .C(n2865), .Y(n3984) );
  NAND2X1 U1064 ( .A(arr[507]), .B(n1259), .Y(n2865) );
  OAI21X1 U1065 ( .A(n2315), .B(n1258), .C(n2866), .Y(n3985) );
  NAND2X1 U1066 ( .A(arr[508]), .B(n1259), .Y(n2866) );
  OAI21X1 U1067 ( .A(n2317), .B(n1258), .C(n2867), .Y(n3986) );
  NAND2X1 U1068 ( .A(arr[509]), .B(n1259), .Y(n2867) );
  OAI21X1 U1069 ( .A(n2319), .B(n1258), .C(n2868), .Y(n3987) );
  NAND2X1 U1070 ( .A(arr[510]), .B(n1259), .Y(n2868) );
  OAI21X1 U1071 ( .A(n2321), .B(n1258), .C(n2869), .Y(n3988) );
  NAND2X1 U1072 ( .A(arr[511]), .B(n1259), .Y(n2869) );
  AND2X1 U1075 ( .A(n2870), .B(n2871), .Y(n2851) );
  OAI21X1 U1076 ( .A(n2291), .B(n1256), .C(n2873), .Y(n3989) );
  NAND2X1 U1077 ( .A(arr[512]), .B(n1257), .Y(n2873) );
  OAI21X1 U1078 ( .A(n2293), .B(n1256), .C(n2874), .Y(n3990) );
  NAND2X1 U1079 ( .A(arr[513]), .B(n1257), .Y(n2874) );
  OAI21X1 U1080 ( .A(n2295), .B(n1256), .C(n2875), .Y(n3991) );
  NAND2X1 U1081 ( .A(arr[514]), .B(n1256), .Y(n2875) );
  OAI21X1 U1082 ( .A(n2297), .B(n1256), .C(n2876), .Y(n3992) );
  NAND2X1 U1083 ( .A(arr[515]), .B(n1256), .Y(n2876) );
  OAI21X1 U1084 ( .A(n2299), .B(n1256), .C(n2877), .Y(n3993) );
  NAND2X1 U1085 ( .A(arr[516]), .B(n1257), .Y(n2877) );
  OAI21X1 U1086 ( .A(n2301), .B(n1256), .C(n2878), .Y(n3994) );
  NAND2X1 U1087 ( .A(arr[517]), .B(n1257), .Y(n2878) );
  OAI21X1 U1088 ( .A(n2303), .B(n1256), .C(n2879), .Y(n3995) );
  NAND2X1 U1089 ( .A(arr[518]), .B(n1257), .Y(n2879) );
  OAI21X1 U1090 ( .A(n2305), .B(n1256), .C(n2880), .Y(n3996) );
  NAND2X1 U1091 ( .A(arr[519]), .B(n1257), .Y(n2880) );
  OAI21X1 U1092 ( .A(n2307), .B(n1256), .C(n2881), .Y(n3997) );
  NAND2X1 U1093 ( .A(arr[520]), .B(n1257), .Y(n2881) );
  OAI21X1 U1094 ( .A(n2309), .B(n1257), .C(n2882), .Y(n3998) );
  NAND2X1 U1095 ( .A(arr[521]), .B(n1257), .Y(n2882) );
  OAI21X1 U1096 ( .A(n2311), .B(n1257), .C(n2883), .Y(n3999) );
  NAND2X1 U1097 ( .A(arr[522]), .B(n1257), .Y(n2883) );
  OAI21X1 U1098 ( .A(n2313), .B(n1257), .C(n2884), .Y(n4000) );
  NAND2X1 U1099 ( .A(arr[523]), .B(n1257), .Y(n2884) );
  OAI21X1 U1100 ( .A(n2315), .B(n1256), .C(n2885), .Y(n4001) );
  NAND2X1 U1101 ( .A(arr[524]), .B(n1257), .Y(n2885) );
  OAI21X1 U1102 ( .A(n2317), .B(n1256), .C(n2886), .Y(n4002) );
  NAND2X1 U1103 ( .A(arr[525]), .B(n1257), .Y(n2886) );
  OAI21X1 U1104 ( .A(n2319), .B(n1256), .C(n2887), .Y(n4003) );
  NAND2X1 U1105 ( .A(arr[526]), .B(n1257), .Y(n2887) );
  OAI21X1 U1106 ( .A(n2321), .B(n1256), .C(n2888), .Y(n4004) );
  NAND2X1 U1107 ( .A(arr[527]), .B(n1257), .Y(n2888) );
  OAI21X1 U1109 ( .A(n2291), .B(n1254), .C(n2891), .Y(n4005) );
  NAND2X1 U1110 ( .A(arr[528]), .B(n1255), .Y(n2891) );
  OAI21X1 U1111 ( .A(n2293), .B(n1254), .C(n2892), .Y(n4006) );
  NAND2X1 U1112 ( .A(arr[529]), .B(n1255), .Y(n2892) );
  OAI21X1 U1113 ( .A(n2295), .B(n1254), .C(n2893), .Y(n4007) );
  NAND2X1 U1114 ( .A(arr[530]), .B(n1254), .Y(n2893) );
  OAI21X1 U1115 ( .A(n2297), .B(n1254), .C(n2894), .Y(n4008) );
  NAND2X1 U1116 ( .A(arr[531]), .B(n1254), .Y(n2894) );
  OAI21X1 U1117 ( .A(n2299), .B(n1254), .C(n2895), .Y(n4009) );
  NAND2X1 U1118 ( .A(arr[532]), .B(n1255), .Y(n2895) );
  OAI21X1 U1119 ( .A(n2301), .B(n1254), .C(n2896), .Y(n4010) );
  NAND2X1 U1120 ( .A(arr[533]), .B(n1255), .Y(n2896) );
  OAI21X1 U1121 ( .A(n2303), .B(n1254), .C(n2897), .Y(n4011) );
  NAND2X1 U1122 ( .A(arr[534]), .B(n1255), .Y(n2897) );
  OAI21X1 U1123 ( .A(n2305), .B(n1254), .C(n2898), .Y(n4012) );
  NAND2X1 U1124 ( .A(arr[535]), .B(n1255), .Y(n2898) );
  OAI21X1 U1125 ( .A(n2307), .B(n1254), .C(n2899), .Y(n4013) );
  NAND2X1 U1126 ( .A(arr[536]), .B(n1255), .Y(n2899) );
  OAI21X1 U1127 ( .A(n2309), .B(n1255), .C(n2900), .Y(n4014) );
  NAND2X1 U1128 ( .A(arr[537]), .B(n1255), .Y(n2900) );
  OAI21X1 U1129 ( .A(n2311), .B(n1255), .C(n2901), .Y(n4015) );
  NAND2X1 U1130 ( .A(arr[538]), .B(n1255), .Y(n2901) );
  OAI21X1 U1131 ( .A(n2313), .B(n1255), .C(n2902), .Y(n4016) );
  NAND2X1 U1132 ( .A(arr[539]), .B(n1255), .Y(n2902) );
  OAI21X1 U1133 ( .A(n2315), .B(n1254), .C(n2903), .Y(n4017) );
  NAND2X1 U1134 ( .A(arr[540]), .B(n1255), .Y(n2903) );
  OAI21X1 U1135 ( .A(n2317), .B(n1254), .C(n2904), .Y(n4018) );
  NAND2X1 U1136 ( .A(arr[541]), .B(n1255), .Y(n2904) );
  OAI21X1 U1137 ( .A(n2319), .B(n1254), .C(n2905), .Y(n4019) );
  NAND2X1 U1138 ( .A(arr[542]), .B(n1255), .Y(n2905) );
  OAI21X1 U1139 ( .A(n2321), .B(n1254), .C(n2906), .Y(n4020) );
  NAND2X1 U1140 ( .A(arr[543]), .B(n1255), .Y(n2906) );
  AND2X1 U1142 ( .A(n2908), .B(n2909), .Y(n2324) );
  OAI21X1 U1143 ( .A(n2291), .B(n1252), .C(n2911), .Y(n4021) );
  NAND2X1 U1144 ( .A(arr[544]), .B(n1253), .Y(n2911) );
  OAI21X1 U1145 ( .A(n2293), .B(n1252), .C(n2912), .Y(n4022) );
  NAND2X1 U1146 ( .A(arr[545]), .B(n1253), .Y(n2912) );
  OAI21X1 U1147 ( .A(n2295), .B(n1252), .C(n2913), .Y(n4023) );
  NAND2X1 U1148 ( .A(arr[546]), .B(n1252), .Y(n2913) );
  OAI21X1 U1149 ( .A(n2297), .B(n1252), .C(n2914), .Y(n4024) );
  NAND2X1 U1150 ( .A(arr[547]), .B(n1252), .Y(n2914) );
  OAI21X1 U1151 ( .A(n2299), .B(n1252), .C(n2915), .Y(n4025) );
  NAND2X1 U1152 ( .A(arr[548]), .B(n1253), .Y(n2915) );
  OAI21X1 U1153 ( .A(n2301), .B(n1252), .C(n2916), .Y(n4026) );
  NAND2X1 U1154 ( .A(arr[549]), .B(n1253), .Y(n2916) );
  OAI21X1 U1155 ( .A(n2303), .B(n1252), .C(n2917), .Y(n4027) );
  NAND2X1 U1156 ( .A(arr[550]), .B(n1253), .Y(n2917) );
  OAI21X1 U1157 ( .A(n2305), .B(n1252), .C(n2918), .Y(n4028) );
  NAND2X1 U1158 ( .A(arr[551]), .B(n1253), .Y(n2918) );
  OAI21X1 U1159 ( .A(n2307), .B(n1252), .C(n2919), .Y(n4029) );
  NAND2X1 U1160 ( .A(arr[552]), .B(n1253), .Y(n2919) );
  OAI21X1 U1161 ( .A(n2309), .B(n1253), .C(n2920), .Y(n4030) );
  NAND2X1 U1162 ( .A(arr[553]), .B(n1253), .Y(n2920) );
  OAI21X1 U1163 ( .A(n2311), .B(n1253), .C(n2921), .Y(n4031) );
  NAND2X1 U1164 ( .A(arr[554]), .B(n1253), .Y(n2921) );
  OAI21X1 U1165 ( .A(n2313), .B(n1253), .C(n2922), .Y(n4032) );
  NAND2X1 U1166 ( .A(arr[555]), .B(n1253), .Y(n2922) );
  OAI21X1 U1167 ( .A(n2315), .B(n1252), .C(n2923), .Y(n4033) );
  NAND2X1 U1168 ( .A(arr[556]), .B(n1253), .Y(n2923) );
  OAI21X1 U1169 ( .A(n2317), .B(n1252), .C(n2924), .Y(n4034) );
  NAND2X1 U1170 ( .A(arr[557]), .B(n1253), .Y(n2924) );
  OAI21X1 U1171 ( .A(n2319), .B(n1252), .C(n2925), .Y(n4035) );
  NAND2X1 U1172 ( .A(arr[558]), .B(n1253), .Y(n2925) );
  OAI21X1 U1173 ( .A(n2321), .B(n1252), .C(n2926), .Y(n4036) );
  NAND2X1 U1174 ( .A(arr[559]), .B(n1253), .Y(n2926) );
  OAI21X1 U1176 ( .A(n2291), .B(n1250), .C(n2928), .Y(n4037) );
  NAND2X1 U1177 ( .A(arr[560]), .B(n1251), .Y(n2928) );
  OAI21X1 U1178 ( .A(n2293), .B(n1250), .C(n2929), .Y(n4038) );
  NAND2X1 U1179 ( .A(arr[561]), .B(n1251), .Y(n2929) );
  OAI21X1 U1180 ( .A(n2295), .B(n1250), .C(n2930), .Y(n4039) );
  NAND2X1 U1181 ( .A(arr[562]), .B(n1250), .Y(n2930) );
  OAI21X1 U1182 ( .A(n2297), .B(n1250), .C(n2931), .Y(n4040) );
  NAND2X1 U1183 ( .A(arr[563]), .B(n1250), .Y(n2931) );
  OAI21X1 U1184 ( .A(n2299), .B(n1250), .C(n2932), .Y(n4041) );
  NAND2X1 U1185 ( .A(arr[564]), .B(n1251), .Y(n2932) );
  OAI21X1 U1186 ( .A(n2301), .B(n1250), .C(n2933), .Y(n4042) );
  NAND2X1 U1187 ( .A(arr[565]), .B(n1251), .Y(n2933) );
  OAI21X1 U1188 ( .A(n2303), .B(n1250), .C(n2934), .Y(n4043) );
  NAND2X1 U1189 ( .A(arr[566]), .B(n1251), .Y(n2934) );
  OAI21X1 U1190 ( .A(n2305), .B(n1250), .C(n2935), .Y(n4044) );
  NAND2X1 U1191 ( .A(arr[567]), .B(n1251), .Y(n2935) );
  OAI21X1 U1192 ( .A(n2307), .B(n1250), .C(n2936), .Y(n4045) );
  NAND2X1 U1193 ( .A(arr[568]), .B(n1251), .Y(n2936) );
  OAI21X1 U1194 ( .A(n2309), .B(n1251), .C(n2937), .Y(n4046) );
  NAND2X1 U1195 ( .A(arr[569]), .B(n1251), .Y(n2937) );
  OAI21X1 U1196 ( .A(n2311), .B(n1251), .C(n2938), .Y(n4047) );
  NAND2X1 U1197 ( .A(arr[570]), .B(n1251), .Y(n2938) );
  OAI21X1 U1198 ( .A(n2313), .B(n1251), .C(n2939), .Y(n4048) );
  NAND2X1 U1199 ( .A(arr[571]), .B(n1251), .Y(n2939) );
  OAI21X1 U1200 ( .A(n2315), .B(n1250), .C(n2940), .Y(n4049) );
  NAND2X1 U1201 ( .A(arr[572]), .B(n1251), .Y(n2940) );
  OAI21X1 U1202 ( .A(n2317), .B(n1250), .C(n2941), .Y(n4050) );
  NAND2X1 U1203 ( .A(arr[573]), .B(n1251), .Y(n2941) );
  OAI21X1 U1204 ( .A(n2319), .B(n1250), .C(n2942), .Y(n4051) );
  NAND2X1 U1205 ( .A(arr[574]), .B(n1251), .Y(n2942) );
  OAI21X1 U1206 ( .A(n2321), .B(n1250), .C(n2943), .Y(n4052) );
  NAND2X1 U1207 ( .A(arr[575]), .B(n1251), .Y(n2943) );
  AND2X1 U1209 ( .A(n2944), .B(n2908), .Y(n2360) );
  OAI21X1 U1210 ( .A(n2291), .B(n1248), .C(n2946), .Y(n4053) );
  NAND2X1 U1211 ( .A(arr[576]), .B(n1249), .Y(n2946) );
  OAI21X1 U1212 ( .A(n2293), .B(n1248), .C(n2947), .Y(n4054) );
  NAND2X1 U1213 ( .A(arr[577]), .B(n1249), .Y(n2947) );
  OAI21X1 U1214 ( .A(n2295), .B(n1248), .C(n2948), .Y(n4055) );
  NAND2X1 U1215 ( .A(arr[578]), .B(n1248), .Y(n2948) );
  OAI21X1 U1216 ( .A(n2297), .B(n1248), .C(n2949), .Y(n4056) );
  NAND2X1 U1217 ( .A(arr[579]), .B(n1248), .Y(n2949) );
  OAI21X1 U1218 ( .A(n2299), .B(n1248), .C(n2950), .Y(n4057) );
  NAND2X1 U1219 ( .A(arr[580]), .B(n1249), .Y(n2950) );
  OAI21X1 U1220 ( .A(n2301), .B(n1248), .C(n2951), .Y(n4058) );
  NAND2X1 U1221 ( .A(arr[581]), .B(n1249), .Y(n2951) );
  OAI21X1 U1222 ( .A(n2303), .B(n1248), .C(n2952), .Y(n4059) );
  NAND2X1 U1223 ( .A(arr[582]), .B(n1249), .Y(n2952) );
  OAI21X1 U1224 ( .A(n2305), .B(n1248), .C(n2953), .Y(n4060) );
  NAND2X1 U1225 ( .A(arr[583]), .B(n1249), .Y(n2953) );
  OAI21X1 U1226 ( .A(n2307), .B(n1248), .C(n2954), .Y(n4061) );
  NAND2X1 U1227 ( .A(arr[584]), .B(n1249), .Y(n2954) );
  OAI21X1 U1228 ( .A(n2309), .B(n1249), .C(n2955), .Y(n4062) );
  NAND2X1 U1229 ( .A(arr[585]), .B(n1249), .Y(n2955) );
  OAI21X1 U1230 ( .A(n2311), .B(n1249), .C(n2956), .Y(n4063) );
  NAND2X1 U1231 ( .A(arr[586]), .B(n1249), .Y(n2956) );
  OAI21X1 U1232 ( .A(n2313), .B(n1249), .C(n2957), .Y(n4064) );
  NAND2X1 U1233 ( .A(arr[587]), .B(n1249), .Y(n2957) );
  OAI21X1 U1234 ( .A(n2315), .B(n1248), .C(n2958), .Y(n4065) );
  NAND2X1 U1235 ( .A(arr[588]), .B(n1249), .Y(n2958) );
  OAI21X1 U1236 ( .A(n2317), .B(n1248), .C(n2959), .Y(n4066) );
  NAND2X1 U1237 ( .A(arr[589]), .B(n1249), .Y(n2959) );
  OAI21X1 U1238 ( .A(n2319), .B(n1248), .C(n2960), .Y(n4067) );
  NAND2X1 U1239 ( .A(arr[590]), .B(n1249), .Y(n2960) );
  OAI21X1 U1240 ( .A(n2321), .B(n1248), .C(n2961), .Y(n4068) );
  NAND2X1 U1241 ( .A(arr[591]), .B(n1249), .Y(n2961) );
  OAI21X1 U1243 ( .A(n2291), .B(n1246), .C(n2963), .Y(n4069) );
  NAND2X1 U1244 ( .A(arr[592]), .B(n1247), .Y(n2963) );
  OAI21X1 U1245 ( .A(n2293), .B(n1246), .C(n2964), .Y(n4070) );
  NAND2X1 U1246 ( .A(arr[593]), .B(n1247), .Y(n2964) );
  OAI21X1 U1247 ( .A(n2295), .B(n1246), .C(n2965), .Y(n4071) );
  NAND2X1 U1248 ( .A(arr[594]), .B(n1246), .Y(n2965) );
  OAI21X1 U1249 ( .A(n2297), .B(n1246), .C(n2966), .Y(n4072) );
  NAND2X1 U1250 ( .A(arr[595]), .B(n1246), .Y(n2966) );
  OAI21X1 U1251 ( .A(n2299), .B(n1246), .C(n2967), .Y(n4073) );
  NAND2X1 U1252 ( .A(arr[596]), .B(n1247), .Y(n2967) );
  OAI21X1 U1253 ( .A(n2301), .B(n1246), .C(n2968), .Y(n4074) );
  NAND2X1 U1254 ( .A(arr[597]), .B(n1247), .Y(n2968) );
  OAI21X1 U1255 ( .A(n2303), .B(n1246), .C(n2969), .Y(n4075) );
  NAND2X1 U1256 ( .A(arr[598]), .B(n1247), .Y(n2969) );
  OAI21X1 U1257 ( .A(n2305), .B(n1246), .C(n2970), .Y(n4076) );
  NAND2X1 U1258 ( .A(arr[599]), .B(n1247), .Y(n2970) );
  OAI21X1 U1259 ( .A(n2307), .B(n1246), .C(n2971), .Y(n4077) );
  NAND2X1 U1260 ( .A(arr[600]), .B(n1247), .Y(n2971) );
  OAI21X1 U1261 ( .A(n2309), .B(n1247), .C(n2972), .Y(n4078) );
  NAND2X1 U1262 ( .A(arr[601]), .B(n1247), .Y(n2972) );
  OAI21X1 U1263 ( .A(n2311), .B(n1247), .C(n2973), .Y(n4079) );
  NAND2X1 U1264 ( .A(arr[602]), .B(n1247), .Y(n2973) );
  OAI21X1 U1265 ( .A(n2313), .B(n1247), .C(n2974), .Y(n4080) );
  NAND2X1 U1266 ( .A(arr[603]), .B(n1247), .Y(n2974) );
  OAI21X1 U1267 ( .A(n2315), .B(n1246), .C(n2975), .Y(n4081) );
  NAND2X1 U1268 ( .A(arr[604]), .B(n1247), .Y(n2975) );
  OAI21X1 U1269 ( .A(n2317), .B(n1246), .C(n2976), .Y(n4082) );
  NAND2X1 U1270 ( .A(arr[605]), .B(n1247), .Y(n2976) );
  OAI21X1 U1271 ( .A(n2319), .B(n1246), .C(n2977), .Y(n4083) );
  NAND2X1 U1272 ( .A(arr[606]), .B(n1247), .Y(n2977) );
  OAI21X1 U1273 ( .A(n2321), .B(n1246), .C(n2978), .Y(n4084) );
  NAND2X1 U1274 ( .A(arr[607]), .B(n1247), .Y(n2978) );
  AND2X1 U1276 ( .A(n2979), .B(n2908), .Y(n2395) );
  OAI21X1 U1277 ( .A(n2291), .B(n1244), .C(n2981), .Y(n4085) );
  NAND2X1 U1278 ( .A(arr[608]), .B(n1245), .Y(n2981) );
  OAI21X1 U1279 ( .A(n2293), .B(n1244), .C(n2982), .Y(n4086) );
  NAND2X1 U1280 ( .A(arr[609]), .B(n1245), .Y(n2982) );
  OAI21X1 U1281 ( .A(n2295), .B(n1244), .C(n2983), .Y(n4087) );
  NAND2X1 U1282 ( .A(arr[610]), .B(n1244), .Y(n2983) );
  OAI21X1 U1283 ( .A(n2297), .B(n1244), .C(n2984), .Y(n4088) );
  NAND2X1 U1284 ( .A(arr[611]), .B(n1244), .Y(n2984) );
  OAI21X1 U1285 ( .A(n2299), .B(n1244), .C(n2985), .Y(n4089) );
  NAND2X1 U1286 ( .A(arr[612]), .B(n1245), .Y(n2985) );
  OAI21X1 U1287 ( .A(n2301), .B(n1244), .C(n2986), .Y(n4090) );
  NAND2X1 U1288 ( .A(arr[613]), .B(n1245), .Y(n2986) );
  OAI21X1 U1289 ( .A(n2303), .B(n1244), .C(n2987), .Y(n4091) );
  NAND2X1 U1290 ( .A(arr[614]), .B(n1245), .Y(n2987) );
  OAI21X1 U1291 ( .A(n2305), .B(n1244), .C(n2988), .Y(n4092) );
  NAND2X1 U1292 ( .A(arr[615]), .B(n1245), .Y(n2988) );
  OAI21X1 U1293 ( .A(n2307), .B(n1244), .C(n2989), .Y(n4093) );
  NAND2X1 U1294 ( .A(arr[616]), .B(n1245), .Y(n2989) );
  OAI21X1 U1295 ( .A(n2309), .B(n1245), .C(n2990), .Y(n4094) );
  NAND2X1 U1296 ( .A(arr[617]), .B(n1245), .Y(n2990) );
  OAI21X1 U1297 ( .A(n2311), .B(n1245), .C(n2991), .Y(n4095) );
  NAND2X1 U1298 ( .A(arr[618]), .B(n1245), .Y(n2991) );
  OAI21X1 U1299 ( .A(n2313), .B(n1245), .C(n2992), .Y(n4096) );
  NAND2X1 U1300 ( .A(arr[619]), .B(n1245), .Y(n2992) );
  OAI21X1 U1301 ( .A(n2315), .B(n1244), .C(n2993), .Y(n4097) );
  NAND2X1 U1302 ( .A(arr[620]), .B(n1245), .Y(n2993) );
  OAI21X1 U1303 ( .A(n2317), .B(n1244), .C(n2994), .Y(n4098) );
  NAND2X1 U1304 ( .A(arr[621]), .B(n1245), .Y(n2994) );
  OAI21X1 U1305 ( .A(n2319), .B(n1244), .C(n2995), .Y(n4099) );
  NAND2X1 U1306 ( .A(arr[622]), .B(n1245), .Y(n2995) );
  OAI21X1 U1307 ( .A(n2321), .B(n1244), .C(n2996), .Y(n4100) );
  NAND2X1 U1308 ( .A(arr[623]), .B(n1245), .Y(n2996) );
  OAI21X1 U1310 ( .A(n1335), .B(n1242), .C(n2998), .Y(n4101) );
  NAND2X1 U1311 ( .A(arr[624]), .B(n1243), .Y(n2998) );
  OAI21X1 U1312 ( .A(n1334), .B(n1242), .C(n2999), .Y(n4102) );
  NAND2X1 U1313 ( .A(arr[625]), .B(n1243), .Y(n2999) );
  OAI21X1 U1314 ( .A(n1333), .B(n1242), .C(n3000), .Y(n4103) );
  NAND2X1 U1315 ( .A(arr[626]), .B(n1242), .Y(n3000) );
  OAI21X1 U1316 ( .A(n1332), .B(n1242), .C(n3001), .Y(n4104) );
  NAND2X1 U1317 ( .A(arr[627]), .B(n1242), .Y(n3001) );
  OAI21X1 U1318 ( .A(n1331), .B(n1242), .C(n3002), .Y(n4105) );
  NAND2X1 U1319 ( .A(arr[628]), .B(n1243), .Y(n3002) );
  OAI21X1 U1320 ( .A(n1330), .B(n1242), .C(n3003), .Y(n4106) );
  NAND2X1 U1321 ( .A(arr[629]), .B(n1243), .Y(n3003) );
  OAI21X1 U1322 ( .A(n1329), .B(n1242), .C(n3004), .Y(n4107) );
  NAND2X1 U1323 ( .A(arr[630]), .B(n1243), .Y(n3004) );
  OAI21X1 U1324 ( .A(n1328), .B(n1242), .C(n3005), .Y(n4108) );
  NAND2X1 U1325 ( .A(arr[631]), .B(n1243), .Y(n3005) );
  OAI21X1 U1326 ( .A(n1327), .B(n1242), .C(n3006), .Y(n4109) );
  NAND2X1 U1327 ( .A(arr[632]), .B(n1243), .Y(n3006) );
  OAI21X1 U1328 ( .A(n1326), .B(n1243), .C(n3007), .Y(n4110) );
  NAND2X1 U1329 ( .A(arr[633]), .B(n1243), .Y(n3007) );
  OAI21X1 U1330 ( .A(n1325), .B(n1243), .C(n3008), .Y(n4111) );
  NAND2X1 U1331 ( .A(arr[634]), .B(n1243), .Y(n3008) );
  OAI21X1 U1332 ( .A(n1324), .B(n1243), .C(n3009), .Y(n4112) );
  NAND2X1 U1333 ( .A(arr[635]), .B(n1243), .Y(n3009) );
  OAI21X1 U1334 ( .A(n1323), .B(n1242), .C(n3010), .Y(n4113) );
  NAND2X1 U1335 ( .A(arr[636]), .B(n1243), .Y(n3010) );
  OAI21X1 U1336 ( .A(n1322), .B(n1242), .C(n3011), .Y(n4114) );
  NAND2X1 U1337 ( .A(arr[637]), .B(n1243), .Y(n3011) );
  OAI21X1 U1338 ( .A(n1321), .B(n1242), .C(n3012), .Y(n4115) );
  NAND2X1 U1339 ( .A(arr[638]), .B(n1243), .Y(n3012) );
  OAI21X1 U1340 ( .A(n1320), .B(n1242), .C(n3013), .Y(n4116) );
  NAND2X1 U1341 ( .A(arr[639]), .B(n1243), .Y(n3013) );
  AND2X1 U1343 ( .A(n3014), .B(n2908), .Y(n2430) );
  NOR2X1 U1344 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .Y(n2908) );
  OAI21X1 U1345 ( .A(n2291), .B(n1240), .C(n3016), .Y(n4117) );
  NAND2X1 U1346 ( .A(arr[640]), .B(n1241), .Y(n3016) );
  OAI21X1 U1347 ( .A(n2293), .B(n1240), .C(n3017), .Y(n4118) );
  NAND2X1 U1348 ( .A(arr[641]), .B(n1241), .Y(n3017) );
  OAI21X1 U1349 ( .A(n2295), .B(n1240), .C(n3018), .Y(n4119) );
  NAND2X1 U1350 ( .A(arr[642]), .B(n1240), .Y(n3018) );
  OAI21X1 U1351 ( .A(n2297), .B(n1240), .C(n3019), .Y(n4120) );
  NAND2X1 U1352 ( .A(arr[643]), .B(n1240), .Y(n3019) );
  OAI21X1 U1353 ( .A(n2299), .B(n1240), .C(n3020), .Y(n4121) );
  NAND2X1 U1354 ( .A(arr[644]), .B(n1241), .Y(n3020) );
  OAI21X1 U1355 ( .A(n2301), .B(n1240), .C(n3021), .Y(n4122) );
  NAND2X1 U1356 ( .A(arr[645]), .B(n1241), .Y(n3021) );
  OAI21X1 U1357 ( .A(n2303), .B(n1240), .C(n3022), .Y(n4123) );
  NAND2X1 U1358 ( .A(arr[646]), .B(n1241), .Y(n3022) );
  OAI21X1 U1359 ( .A(n2305), .B(n1240), .C(n3023), .Y(n4124) );
  NAND2X1 U1360 ( .A(arr[647]), .B(n1241), .Y(n3023) );
  OAI21X1 U1361 ( .A(n2307), .B(n1240), .C(n3024), .Y(n4125) );
  NAND2X1 U1362 ( .A(arr[648]), .B(n1241), .Y(n3024) );
  OAI21X1 U1363 ( .A(n2309), .B(n1241), .C(n3025), .Y(n4126) );
  NAND2X1 U1364 ( .A(arr[649]), .B(n1241), .Y(n3025) );
  OAI21X1 U1365 ( .A(n2311), .B(n1241), .C(n3026), .Y(n4127) );
  NAND2X1 U1366 ( .A(arr[650]), .B(n1241), .Y(n3026) );
  OAI21X1 U1367 ( .A(n2313), .B(n1241), .C(n3027), .Y(n4128) );
  NAND2X1 U1368 ( .A(arr[651]), .B(n1241), .Y(n3027) );
  OAI21X1 U1369 ( .A(n2315), .B(n1240), .C(n3028), .Y(n4129) );
  NAND2X1 U1370 ( .A(arr[652]), .B(n1241), .Y(n3028) );
  OAI21X1 U1371 ( .A(n2317), .B(n1240), .C(n3029), .Y(n4130) );
  NAND2X1 U1372 ( .A(arr[653]), .B(n1241), .Y(n3029) );
  OAI21X1 U1373 ( .A(n2319), .B(n1240), .C(n3030), .Y(n4131) );
  NAND2X1 U1374 ( .A(arr[654]), .B(n1241), .Y(n3030) );
  OAI21X1 U1375 ( .A(n2321), .B(n1240), .C(n3031), .Y(n4132) );
  NAND2X1 U1376 ( .A(arr[655]), .B(n1241), .Y(n3031) );
  OAI21X1 U1378 ( .A(n2291), .B(n1238), .C(n3033), .Y(n4133) );
  NAND2X1 U1379 ( .A(arr[656]), .B(n1239), .Y(n3033) );
  OAI21X1 U1380 ( .A(n2293), .B(n1238), .C(n3034), .Y(n4134) );
  NAND2X1 U1381 ( .A(arr[657]), .B(n1239), .Y(n3034) );
  OAI21X1 U1382 ( .A(n2295), .B(n1238), .C(n3035), .Y(n4135) );
  NAND2X1 U1383 ( .A(arr[658]), .B(n1238), .Y(n3035) );
  OAI21X1 U1384 ( .A(n2297), .B(n1238), .C(n3036), .Y(n4136) );
  NAND2X1 U1385 ( .A(arr[659]), .B(n1238), .Y(n3036) );
  OAI21X1 U1386 ( .A(n2299), .B(n1238), .C(n3037), .Y(n4137) );
  NAND2X1 U1387 ( .A(arr[660]), .B(n1239), .Y(n3037) );
  OAI21X1 U1388 ( .A(n2301), .B(n1238), .C(n3038), .Y(n4138) );
  NAND2X1 U1389 ( .A(arr[661]), .B(n1239), .Y(n3038) );
  OAI21X1 U1390 ( .A(n2303), .B(n1238), .C(n3039), .Y(n4139) );
  NAND2X1 U1391 ( .A(arr[662]), .B(n1239), .Y(n3039) );
  OAI21X1 U1392 ( .A(n2305), .B(n1238), .C(n3040), .Y(n4140) );
  NAND2X1 U1393 ( .A(arr[663]), .B(n1239), .Y(n3040) );
  OAI21X1 U1394 ( .A(n2307), .B(n1238), .C(n3041), .Y(n4141) );
  NAND2X1 U1395 ( .A(arr[664]), .B(n1239), .Y(n3041) );
  OAI21X1 U1396 ( .A(n2309), .B(n1239), .C(n3042), .Y(n4142) );
  NAND2X1 U1397 ( .A(arr[665]), .B(n1239), .Y(n3042) );
  OAI21X1 U1398 ( .A(n2311), .B(n1239), .C(n3043), .Y(n4143) );
  NAND2X1 U1399 ( .A(arr[666]), .B(n1239), .Y(n3043) );
  OAI21X1 U1400 ( .A(n2313), .B(n1239), .C(n3044), .Y(n4144) );
  NAND2X1 U1401 ( .A(arr[667]), .B(n1239), .Y(n3044) );
  OAI21X1 U1402 ( .A(n2315), .B(n1238), .C(n3045), .Y(n4145) );
  NAND2X1 U1403 ( .A(arr[668]), .B(n1239), .Y(n3045) );
  OAI21X1 U1404 ( .A(n2317), .B(n1238), .C(n3046), .Y(n4146) );
  NAND2X1 U1405 ( .A(arr[669]), .B(n1239), .Y(n3046) );
  OAI21X1 U1406 ( .A(n2319), .B(n1238), .C(n3047), .Y(n4147) );
  NAND2X1 U1407 ( .A(arr[670]), .B(n1239), .Y(n3047) );
  OAI21X1 U1408 ( .A(n2321), .B(n1238), .C(n3048), .Y(n4148) );
  NAND2X1 U1409 ( .A(arr[671]), .B(n1239), .Y(n3048) );
  AND2X1 U1411 ( .A(n3049), .B(n2909), .Y(n2465) );
  OAI21X1 U1412 ( .A(n2291), .B(n1236), .C(n3051), .Y(n4149) );
  NAND2X1 U1413 ( .A(arr[672]), .B(n1237), .Y(n3051) );
  OAI21X1 U1414 ( .A(n2293), .B(n1236), .C(n3052), .Y(n4150) );
  NAND2X1 U1415 ( .A(arr[673]), .B(n1237), .Y(n3052) );
  OAI21X1 U1416 ( .A(n2295), .B(n1236), .C(n3053), .Y(n4151) );
  NAND2X1 U1417 ( .A(arr[674]), .B(n1236), .Y(n3053) );
  OAI21X1 U1418 ( .A(n2297), .B(n1236), .C(n3054), .Y(n4152) );
  NAND2X1 U1419 ( .A(arr[675]), .B(n1236), .Y(n3054) );
  OAI21X1 U1420 ( .A(n2299), .B(n1236), .C(n3055), .Y(n4153) );
  NAND2X1 U1421 ( .A(arr[676]), .B(n1237), .Y(n3055) );
  OAI21X1 U1422 ( .A(n2301), .B(n1236), .C(n3056), .Y(n4154) );
  NAND2X1 U1423 ( .A(arr[677]), .B(n1237), .Y(n3056) );
  OAI21X1 U1424 ( .A(n2303), .B(n1236), .C(n3057), .Y(n4155) );
  NAND2X1 U1425 ( .A(arr[678]), .B(n1237), .Y(n3057) );
  OAI21X1 U1426 ( .A(n2305), .B(n1236), .C(n3058), .Y(n4156) );
  NAND2X1 U1427 ( .A(arr[679]), .B(n1237), .Y(n3058) );
  OAI21X1 U1428 ( .A(n2307), .B(n1236), .C(n3059), .Y(n4157) );
  NAND2X1 U1429 ( .A(arr[680]), .B(n1237), .Y(n3059) );
  OAI21X1 U1430 ( .A(n2309), .B(n1237), .C(n3060), .Y(n4158) );
  NAND2X1 U1431 ( .A(arr[681]), .B(n1237), .Y(n3060) );
  OAI21X1 U1432 ( .A(n2311), .B(n1237), .C(n3061), .Y(n4159) );
  NAND2X1 U1433 ( .A(arr[682]), .B(n1237), .Y(n3061) );
  OAI21X1 U1434 ( .A(n2313), .B(n1237), .C(n3062), .Y(n4160) );
  NAND2X1 U1435 ( .A(arr[683]), .B(n1237), .Y(n3062) );
  OAI21X1 U1436 ( .A(n2315), .B(n1236), .C(n3063), .Y(n4161) );
  NAND2X1 U1437 ( .A(arr[684]), .B(n1237), .Y(n3063) );
  OAI21X1 U1438 ( .A(n2317), .B(n1236), .C(n3064), .Y(n4162) );
  NAND2X1 U1439 ( .A(arr[685]), .B(n1237), .Y(n3064) );
  OAI21X1 U1440 ( .A(n2319), .B(n1236), .C(n3065), .Y(n4163) );
  NAND2X1 U1441 ( .A(arr[686]), .B(n1237), .Y(n3065) );
  OAI21X1 U1442 ( .A(n2321), .B(n1236), .C(n3066), .Y(n4164) );
  NAND2X1 U1443 ( .A(arr[687]), .B(n1237), .Y(n3066) );
  OAI21X1 U1445 ( .A(n1335), .B(n1234), .C(n3068), .Y(n4165) );
  NAND2X1 U1446 ( .A(arr[688]), .B(n1235), .Y(n3068) );
  OAI21X1 U1447 ( .A(n1334), .B(n1234), .C(n3069), .Y(n4166) );
  NAND2X1 U1448 ( .A(arr[689]), .B(n1235), .Y(n3069) );
  OAI21X1 U1449 ( .A(n1333), .B(n1234), .C(n3070), .Y(n4167) );
  NAND2X1 U1450 ( .A(arr[690]), .B(n1234), .Y(n3070) );
  OAI21X1 U1451 ( .A(n1332), .B(n1234), .C(n3071), .Y(n4168) );
  NAND2X1 U1452 ( .A(arr[691]), .B(n1234), .Y(n3071) );
  OAI21X1 U1453 ( .A(n1331), .B(n1234), .C(n3072), .Y(n4169) );
  NAND2X1 U1454 ( .A(arr[692]), .B(n1235), .Y(n3072) );
  OAI21X1 U1455 ( .A(n1330), .B(n1234), .C(n3073), .Y(n4170) );
  NAND2X1 U1456 ( .A(arr[693]), .B(n1235), .Y(n3073) );
  OAI21X1 U1457 ( .A(n1329), .B(n1234), .C(n3074), .Y(n4171) );
  NAND2X1 U1458 ( .A(arr[694]), .B(n1235), .Y(n3074) );
  OAI21X1 U1459 ( .A(n1328), .B(n1234), .C(n3075), .Y(n4172) );
  NAND2X1 U1460 ( .A(arr[695]), .B(n1235), .Y(n3075) );
  OAI21X1 U1461 ( .A(n1327), .B(n1234), .C(n3076), .Y(n4173) );
  NAND2X1 U1462 ( .A(arr[696]), .B(n1235), .Y(n3076) );
  OAI21X1 U1463 ( .A(n1326), .B(n1235), .C(n3077), .Y(n4174) );
  NAND2X1 U1464 ( .A(arr[697]), .B(n1235), .Y(n3077) );
  OAI21X1 U1465 ( .A(n1325), .B(n1235), .C(n3078), .Y(n4175) );
  NAND2X1 U1466 ( .A(arr[698]), .B(n1235), .Y(n3078) );
  OAI21X1 U1467 ( .A(n1324), .B(n1235), .C(n3079), .Y(n4176) );
  NAND2X1 U1468 ( .A(arr[699]), .B(n1235), .Y(n3079) );
  OAI21X1 U1469 ( .A(n1323), .B(n1234), .C(n3080), .Y(n4177) );
  NAND2X1 U1470 ( .A(arr[700]), .B(n1235), .Y(n3080) );
  OAI21X1 U1471 ( .A(n1322), .B(n1234), .C(n3081), .Y(n4178) );
  NAND2X1 U1472 ( .A(arr[701]), .B(n1235), .Y(n3081) );
  OAI21X1 U1473 ( .A(n1321), .B(n1234), .C(n3082), .Y(n4179) );
  NAND2X1 U1474 ( .A(arr[702]), .B(n1235), .Y(n3082) );
  OAI21X1 U1475 ( .A(n1320), .B(n1234), .C(n3083), .Y(n4180) );
  NAND2X1 U1476 ( .A(arr[703]), .B(n1235), .Y(n3083) );
  AND2X1 U1478 ( .A(n3049), .B(n2944), .Y(n2500) );
  OAI21X1 U1479 ( .A(n2291), .B(n1232), .C(n3085), .Y(n4181) );
  NAND2X1 U1480 ( .A(arr[704]), .B(n1233), .Y(n3085) );
  OAI21X1 U1481 ( .A(n2293), .B(n1232), .C(n3086), .Y(n4182) );
  NAND2X1 U1482 ( .A(arr[705]), .B(n1233), .Y(n3086) );
  OAI21X1 U1483 ( .A(n2295), .B(n1232), .C(n3087), .Y(n4183) );
  NAND2X1 U1484 ( .A(arr[706]), .B(n1232), .Y(n3087) );
  OAI21X1 U1485 ( .A(n2297), .B(n1232), .C(n3088), .Y(n4184) );
  NAND2X1 U1486 ( .A(arr[707]), .B(n1232), .Y(n3088) );
  OAI21X1 U1487 ( .A(n2299), .B(n1232), .C(n3089), .Y(n4185) );
  NAND2X1 U1488 ( .A(arr[708]), .B(n1233), .Y(n3089) );
  OAI21X1 U1489 ( .A(n2301), .B(n1232), .C(n3090), .Y(n4186) );
  NAND2X1 U1490 ( .A(arr[709]), .B(n1233), .Y(n3090) );
  OAI21X1 U1491 ( .A(n2303), .B(n1232), .C(n3091), .Y(n4187) );
  NAND2X1 U1492 ( .A(arr[710]), .B(n1233), .Y(n3091) );
  OAI21X1 U1493 ( .A(n2305), .B(n1232), .C(n3092), .Y(n4188) );
  NAND2X1 U1494 ( .A(arr[711]), .B(n1233), .Y(n3092) );
  OAI21X1 U1495 ( .A(n2307), .B(n1232), .C(n3093), .Y(n4189) );
  NAND2X1 U1496 ( .A(arr[712]), .B(n1233), .Y(n3093) );
  OAI21X1 U1497 ( .A(n2309), .B(n1233), .C(n3094), .Y(n4190) );
  NAND2X1 U1498 ( .A(arr[713]), .B(n1233), .Y(n3094) );
  OAI21X1 U1499 ( .A(n2311), .B(n1233), .C(n3095), .Y(n4191) );
  NAND2X1 U1500 ( .A(arr[714]), .B(n1233), .Y(n3095) );
  OAI21X1 U1501 ( .A(n2313), .B(n1233), .C(n3096), .Y(n4192) );
  NAND2X1 U1502 ( .A(arr[715]), .B(n1233), .Y(n3096) );
  OAI21X1 U1503 ( .A(n2315), .B(n1232), .C(n3097), .Y(n4193) );
  NAND2X1 U1504 ( .A(arr[716]), .B(n1233), .Y(n3097) );
  OAI21X1 U1505 ( .A(n2317), .B(n1232), .C(n3098), .Y(n4194) );
  NAND2X1 U1506 ( .A(arr[717]), .B(n1233), .Y(n3098) );
  OAI21X1 U1507 ( .A(n2319), .B(n1232), .C(n3099), .Y(n4195) );
  NAND2X1 U1508 ( .A(arr[718]), .B(n1233), .Y(n3099) );
  OAI21X1 U1509 ( .A(n2321), .B(n1232), .C(n3100), .Y(n4196) );
  NAND2X1 U1510 ( .A(arr[719]), .B(n1233), .Y(n3100) );
  OAI21X1 U1512 ( .A(n2291), .B(n1230), .C(n3102), .Y(n4197) );
  NAND2X1 U1513 ( .A(arr[720]), .B(n1231), .Y(n3102) );
  OAI21X1 U1514 ( .A(n2293), .B(n1230), .C(n3103), .Y(n4198) );
  NAND2X1 U1515 ( .A(arr[721]), .B(n1231), .Y(n3103) );
  OAI21X1 U1516 ( .A(n2295), .B(n1230), .C(n3104), .Y(n4199) );
  NAND2X1 U1517 ( .A(arr[722]), .B(n1230), .Y(n3104) );
  OAI21X1 U1518 ( .A(n2297), .B(n1230), .C(n3105), .Y(n4200) );
  NAND2X1 U1519 ( .A(arr[723]), .B(n1230), .Y(n3105) );
  OAI21X1 U1520 ( .A(n2299), .B(n1230), .C(n3106), .Y(n4201) );
  NAND2X1 U1521 ( .A(arr[724]), .B(n1231), .Y(n3106) );
  OAI21X1 U1522 ( .A(n2301), .B(n1230), .C(n3107), .Y(n4202) );
  NAND2X1 U1523 ( .A(arr[725]), .B(n1231), .Y(n3107) );
  OAI21X1 U1524 ( .A(n2303), .B(n1230), .C(n3108), .Y(n4203) );
  NAND2X1 U1525 ( .A(arr[726]), .B(n1231), .Y(n3108) );
  OAI21X1 U1526 ( .A(n2305), .B(n1230), .C(n3109), .Y(n4204) );
  NAND2X1 U1527 ( .A(arr[727]), .B(n1231), .Y(n3109) );
  OAI21X1 U1528 ( .A(n2307), .B(n1230), .C(n3110), .Y(n4205) );
  NAND2X1 U1529 ( .A(arr[728]), .B(n1231), .Y(n3110) );
  OAI21X1 U1530 ( .A(n2309), .B(n1231), .C(n3111), .Y(n4206) );
  NAND2X1 U1531 ( .A(arr[729]), .B(n1231), .Y(n3111) );
  OAI21X1 U1532 ( .A(n2311), .B(n1231), .C(n3112), .Y(n4207) );
  NAND2X1 U1533 ( .A(arr[730]), .B(n1231), .Y(n3112) );
  OAI21X1 U1534 ( .A(n2313), .B(n1231), .C(n3113), .Y(n4208) );
  NAND2X1 U1535 ( .A(arr[731]), .B(n1231), .Y(n3113) );
  OAI21X1 U1536 ( .A(n2315), .B(n1230), .C(n3114), .Y(n4209) );
  NAND2X1 U1537 ( .A(arr[732]), .B(n1231), .Y(n3114) );
  OAI21X1 U1538 ( .A(n2317), .B(n1230), .C(n3115), .Y(n4210) );
  NAND2X1 U1539 ( .A(arr[733]), .B(n1231), .Y(n3115) );
  OAI21X1 U1540 ( .A(n2319), .B(n1230), .C(n3116), .Y(n4211) );
  NAND2X1 U1541 ( .A(arr[734]), .B(n1231), .Y(n3116) );
  OAI21X1 U1542 ( .A(n2321), .B(n1230), .C(n3117), .Y(n4212) );
  NAND2X1 U1543 ( .A(arr[735]), .B(n1231), .Y(n3117) );
  AND2X1 U1545 ( .A(n3049), .B(n2979), .Y(n2535) );
  OAI21X1 U1546 ( .A(n2291), .B(n1228), .C(n3119), .Y(n4213) );
  NAND2X1 U1547 ( .A(arr[736]), .B(n1229), .Y(n3119) );
  OAI21X1 U1548 ( .A(n2293), .B(n1228), .C(n3120), .Y(n4214) );
  NAND2X1 U1549 ( .A(arr[737]), .B(n1229), .Y(n3120) );
  OAI21X1 U1550 ( .A(n2295), .B(n1228), .C(n3121), .Y(n4215) );
  NAND2X1 U1551 ( .A(arr[738]), .B(n1228), .Y(n3121) );
  OAI21X1 U1552 ( .A(n2297), .B(n1228), .C(n3122), .Y(n4216) );
  NAND2X1 U1553 ( .A(arr[739]), .B(n1228), .Y(n3122) );
  OAI21X1 U1554 ( .A(n2299), .B(n1228), .C(n3123), .Y(n4217) );
  NAND2X1 U1555 ( .A(arr[740]), .B(n1229), .Y(n3123) );
  OAI21X1 U1556 ( .A(n2301), .B(n1228), .C(n3124), .Y(n4218) );
  NAND2X1 U1557 ( .A(arr[741]), .B(n1229), .Y(n3124) );
  OAI21X1 U1558 ( .A(n2303), .B(n1228), .C(n3125), .Y(n4219) );
  NAND2X1 U1559 ( .A(arr[742]), .B(n1229), .Y(n3125) );
  OAI21X1 U1560 ( .A(n2305), .B(n1228), .C(n3126), .Y(n4220) );
  NAND2X1 U1561 ( .A(arr[743]), .B(n1229), .Y(n3126) );
  OAI21X1 U1562 ( .A(n2307), .B(n1228), .C(n3127), .Y(n4221) );
  NAND2X1 U1563 ( .A(arr[744]), .B(n1229), .Y(n3127) );
  OAI21X1 U1564 ( .A(n2309), .B(n1229), .C(n3128), .Y(n4222) );
  NAND2X1 U1565 ( .A(arr[745]), .B(n1229), .Y(n3128) );
  OAI21X1 U1566 ( .A(n2311), .B(n1229), .C(n3129), .Y(n4223) );
  NAND2X1 U1567 ( .A(arr[746]), .B(n1229), .Y(n3129) );
  OAI21X1 U1568 ( .A(n2313), .B(n1229), .C(n3130), .Y(n4224) );
  NAND2X1 U1569 ( .A(arr[747]), .B(n1229), .Y(n3130) );
  OAI21X1 U1570 ( .A(n2315), .B(n1228), .C(n3131), .Y(n4225) );
  NAND2X1 U1571 ( .A(arr[748]), .B(n1229), .Y(n3131) );
  OAI21X1 U1572 ( .A(n2317), .B(n1228), .C(n3132), .Y(n4226) );
  NAND2X1 U1573 ( .A(arr[749]), .B(n1229), .Y(n3132) );
  OAI21X1 U1574 ( .A(n2319), .B(n1228), .C(n3133), .Y(n4227) );
  NAND2X1 U1575 ( .A(arr[750]), .B(n1229), .Y(n3133) );
  OAI21X1 U1576 ( .A(n2321), .B(n1228), .C(n3134), .Y(n4228) );
  NAND2X1 U1577 ( .A(arr[751]), .B(n1229), .Y(n3134) );
  OAI21X1 U1579 ( .A(n1335), .B(n1226), .C(n3136), .Y(n4229) );
  NAND2X1 U1580 ( .A(arr[752]), .B(n1227), .Y(n3136) );
  OAI21X1 U1581 ( .A(n1334), .B(n1226), .C(n3137), .Y(n4230) );
  NAND2X1 U1582 ( .A(arr[753]), .B(n1227), .Y(n3137) );
  OAI21X1 U1583 ( .A(n1333), .B(n1226), .C(n3138), .Y(n4231) );
  NAND2X1 U1584 ( .A(arr[754]), .B(n1226), .Y(n3138) );
  OAI21X1 U1585 ( .A(n1332), .B(n1226), .C(n3139), .Y(n4232) );
  NAND2X1 U1586 ( .A(arr[755]), .B(n1226), .Y(n3139) );
  OAI21X1 U1587 ( .A(n1331), .B(n1226), .C(n3140), .Y(n4233) );
  NAND2X1 U1588 ( .A(arr[756]), .B(n1227), .Y(n3140) );
  OAI21X1 U1589 ( .A(n1330), .B(n1226), .C(n3141), .Y(n4234) );
  NAND2X1 U1590 ( .A(arr[757]), .B(n1227), .Y(n3141) );
  OAI21X1 U1591 ( .A(n1329), .B(n1226), .C(n3142), .Y(n4235) );
  NAND2X1 U1592 ( .A(arr[758]), .B(n1227), .Y(n3142) );
  OAI21X1 U1593 ( .A(n1328), .B(n1226), .C(n3143), .Y(n4236) );
  NAND2X1 U1594 ( .A(arr[759]), .B(n1227), .Y(n3143) );
  OAI21X1 U1595 ( .A(n1327), .B(n1226), .C(n3144), .Y(n4237) );
  NAND2X1 U1596 ( .A(arr[760]), .B(n1227), .Y(n3144) );
  OAI21X1 U1597 ( .A(n1326), .B(n1227), .C(n3145), .Y(n4238) );
  NAND2X1 U1598 ( .A(arr[761]), .B(n1227), .Y(n3145) );
  OAI21X1 U1599 ( .A(n1325), .B(n1227), .C(n3146), .Y(n4239) );
  NAND2X1 U1600 ( .A(arr[762]), .B(n1227), .Y(n3146) );
  OAI21X1 U1601 ( .A(n1324), .B(n1227), .C(n3147), .Y(n4240) );
  NAND2X1 U1602 ( .A(arr[763]), .B(n1227), .Y(n3147) );
  OAI21X1 U1603 ( .A(n1323), .B(n1226), .C(n3148), .Y(n4241) );
  NAND2X1 U1604 ( .A(arr[764]), .B(n1227), .Y(n3148) );
  OAI21X1 U1605 ( .A(n1322), .B(n1226), .C(n3149), .Y(n4242) );
  NAND2X1 U1606 ( .A(arr[765]), .B(n1227), .Y(n3149) );
  OAI21X1 U1607 ( .A(n1321), .B(n1226), .C(n3150), .Y(n4243) );
  NAND2X1 U1608 ( .A(arr[766]), .B(n1227), .Y(n3150) );
  OAI21X1 U1609 ( .A(n1320), .B(n1226), .C(n3151), .Y(n4244) );
  NAND2X1 U1610 ( .A(arr[767]), .B(n1227), .Y(n3151) );
  AND2X1 U1612 ( .A(n3049), .B(n3014), .Y(n2570) );
  NOR2X1 U1613 ( .A(n3152), .B(wr_ptr[4]), .Y(n3049) );
  OAI21X1 U1614 ( .A(n2291), .B(n1224), .C(n3154), .Y(n4245) );
  NAND2X1 U1615 ( .A(arr[768]), .B(n1225), .Y(n3154) );
  OAI21X1 U1616 ( .A(n2293), .B(n1224), .C(n3155), .Y(n4246) );
  NAND2X1 U1617 ( .A(arr[769]), .B(n1225), .Y(n3155) );
  OAI21X1 U1618 ( .A(n2295), .B(n1224), .C(n3156), .Y(n4247) );
  NAND2X1 U1619 ( .A(arr[770]), .B(n1224), .Y(n3156) );
  OAI21X1 U1620 ( .A(n2297), .B(n1224), .C(n3157), .Y(n4248) );
  NAND2X1 U1621 ( .A(arr[771]), .B(n1224), .Y(n3157) );
  OAI21X1 U1622 ( .A(n2299), .B(n1224), .C(n3158), .Y(n4249) );
  NAND2X1 U1623 ( .A(arr[772]), .B(n1225), .Y(n3158) );
  OAI21X1 U1624 ( .A(n2301), .B(n1224), .C(n3159), .Y(n4250) );
  NAND2X1 U1625 ( .A(arr[773]), .B(n1225), .Y(n3159) );
  OAI21X1 U1626 ( .A(n2303), .B(n1224), .C(n3160), .Y(n4251) );
  NAND2X1 U1627 ( .A(arr[774]), .B(n1225), .Y(n3160) );
  OAI21X1 U1628 ( .A(n2305), .B(n1224), .C(n3161), .Y(n4252) );
  NAND2X1 U1629 ( .A(arr[775]), .B(n1225), .Y(n3161) );
  OAI21X1 U1630 ( .A(n2307), .B(n1224), .C(n3162), .Y(n4253) );
  NAND2X1 U1631 ( .A(arr[776]), .B(n1225), .Y(n3162) );
  OAI21X1 U1632 ( .A(n2309), .B(n1225), .C(n3163), .Y(n4254) );
  NAND2X1 U1633 ( .A(arr[777]), .B(n1225), .Y(n3163) );
  OAI21X1 U1634 ( .A(n2311), .B(n1225), .C(n3164), .Y(n4255) );
  NAND2X1 U1635 ( .A(arr[778]), .B(n1225), .Y(n3164) );
  OAI21X1 U1636 ( .A(n2313), .B(n1225), .C(n3165), .Y(n4256) );
  NAND2X1 U1637 ( .A(arr[779]), .B(n1225), .Y(n3165) );
  OAI21X1 U1638 ( .A(n2315), .B(n1224), .C(n3166), .Y(n4257) );
  NAND2X1 U1639 ( .A(arr[780]), .B(n1225), .Y(n3166) );
  OAI21X1 U1640 ( .A(n2317), .B(n1224), .C(n3167), .Y(n4258) );
  NAND2X1 U1641 ( .A(arr[781]), .B(n1225), .Y(n3167) );
  OAI21X1 U1642 ( .A(n2319), .B(n1224), .C(n3168), .Y(n4259) );
  NAND2X1 U1643 ( .A(arr[782]), .B(n1225), .Y(n3168) );
  OAI21X1 U1644 ( .A(n2321), .B(n1224), .C(n3169), .Y(n4260) );
  NAND2X1 U1645 ( .A(arr[783]), .B(n1225), .Y(n3169) );
  OAI21X1 U1647 ( .A(n2291), .B(n1222), .C(n3171), .Y(n4261) );
  NAND2X1 U1648 ( .A(arr[784]), .B(n1223), .Y(n3171) );
  OAI21X1 U1649 ( .A(n2293), .B(n1222), .C(n3172), .Y(n4262) );
  NAND2X1 U1650 ( .A(arr[785]), .B(n1223), .Y(n3172) );
  OAI21X1 U1651 ( .A(n2295), .B(n1222), .C(n3173), .Y(n4263) );
  NAND2X1 U1652 ( .A(arr[786]), .B(n1222), .Y(n3173) );
  OAI21X1 U1653 ( .A(n2297), .B(n1222), .C(n3174), .Y(n4264) );
  NAND2X1 U1654 ( .A(arr[787]), .B(n1222), .Y(n3174) );
  OAI21X1 U1655 ( .A(n2299), .B(n1222), .C(n3175), .Y(n4265) );
  NAND2X1 U1656 ( .A(arr[788]), .B(n1223), .Y(n3175) );
  OAI21X1 U1657 ( .A(n2301), .B(n1222), .C(n3176), .Y(n4266) );
  NAND2X1 U1658 ( .A(arr[789]), .B(n1223), .Y(n3176) );
  OAI21X1 U1659 ( .A(n2303), .B(n1222), .C(n3177), .Y(n4267) );
  NAND2X1 U1660 ( .A(arr[790]), .B(n1223), .Y(n3177) );
  OAI21X1 U1661 ( .A(n2305), .B(n1222), .C(n3178), .Y(n4268) );
  NAND2X1 U1662 ( .A(arr[791]), .B(n1223), .Y(n3178) );
  OAI21X1 U1663 ( .A(n2307), .B(n1222), .C(n3179), .Y(n4269) );
  NAND2X1 U1664 ( .A(arr[792]), .B(n1223), .Y(n3179) );
  OAI21X1 U1665 ( .A(n2309), .B(n1223), .C(n3180), .Y(n4270) );
  NAND2X1 U1666 ( .A(arr[793]), .B(n1223), .Y(n3180) );
  OAI21X1 U1667 ( .A(n2311), .B(n1223), .C(n3181), .Y(n4271) );
  NAND2X1 U1668 ( .A(arr[794]), .B(n1223), .Y(n3181) );
  OAI21X1 U1669 ( .A(n2313), .B(n1223), .C(n3182), .Y(n4272) );
  NAND2X1 U1670 ( .A(arr[795]), .B(n1223), .Y(n3182) );
  OAI21X1 U1671 ( .A(n2315), .B(n1222), .C(n3183), .Y(n4273) );
  NAND2X1 U1672 ( .A(arr[796]), .B(n1223), .Y(n3183) );
  OAI21X1 U1673 ( .A(n2317), .B(n1222), .C(n3184), .Y(n4274) );
  NAND2X1 U1674 ( .A(arr[797]), .B(n1223), .Y(n3184) );
  OAI21X1 U1675 ( .A(n2319), .B(n1222), .C(n3185), .Y(n4275) );
  NAND2X1 U1676 ( .A(arr[798]), .B(n1223), .Y(n3185) );
  OAI21X1 U1677 ( .A(n2321), .B(n1222), .C(n3186), .Y(n4276) );
  NAND2X1 U1678 ( .A(arr[799]), .B(n1223), .Y(n3186) );
  AND2X1 U1680 ( .A(n3187), .B(n2909), .Y(n2605) );
  OAI21X1 U1681 ( .A(n2291), .B(n1220), .C(n3189), .Y(n4277) );
  NAND2X1 U1682 ( .A(arr[800]), .B(n1221), .Y(n3189) );
  OAI21X1 U1683 ( .A(n2293), .B(n1220), .C(n3190), .Y(n4278) );
  NAND2X1 U1684 ( .A(arr[801]), .B(n1221), .Y(n3190) );
  OAI21X1 U1685 ( .A(n2295), .B(n1220), .C(n3191), .Y(n4279) );
  NAND2X1 U1686 ( .A(arr[802]), .B(n1220), .Y(n3191) );
  OAI21X1 U1687 ( .A(n2297), .B(n1220), .C(n3192), .Y(n4280) );
  NAND2X1 U1688 ( .A(arr[803]), .B(n1220), .Y(n3192) );
  OAI21X1 U1689 ( .A(n2299), .B(n1220), .C(n3193), .Y(n4281) );
  NAND2X1 U1690 ( .A(arr[804]), .B(n1221), .Y(n3193) );
  OAI21X1 U1691 ( .A(n2301), .B(n1220), .C(n3194), .Y(n4282) );
  NAND2X1 U1692 ( .A(arr[805]), .B(n1221), .Y(n3194) );
  OAI21X1 U1693 ( .A(n2303), .B(n1220), .C(n3195), .Y(n4283) );
  NAND2X1 U1694 ( .A(arr[806]), .B(n1221), .Y(n3195) );
  OAI21X1 U1695 ( .A(n2305), .B(n1220), .C(n3196), .Y(n4284) );
  NAND2X1 U1696 ( .A(arr[807]), .B(n1221), .Y(n3196) );
  OAI21X1 U1697 ( .A(n2307), .B(n1220), .C(n3197), .Y(n4285) );
  NAND2X1 U1698 ( .A(arr[808]), .B(n1221), .Y(n3197) );
  OAI21X1 U1699 ( .A(n2309), .B(n1221), .C(n3198), .Y(n4286) );
  NAND2X1 U1700 ( .A(arr[809]), .B(n1221), .Y(n3198) );
  OAI21X1 U1701 ( .A(n2311), .B(n1221), .C(n3199), .Y(n4287) );
  NAND2X1 U1702 ( .A(arr[810]), .B(n1221), .Y(n3199) );
  OAI21X1 U1703 ( .A(n2313), .B(n1221), .C(n3200), .Y(n4288) );
  NAND2X1 U1704 ( .A(arr[811]), .B(n1221), .Y(n3200) );
  OAI21X1 U1705 ( .A(n2315), .B(n1220), .C(n3201), .Y(n4289) );
  NAND2X1 U1706 ( .A(arr[812]), .B(n1221), .Y(n3201) );
  OAI21X1 U1707 ( .A(n2317), .B(n1220), .C(n3202), .Y(n4290) );
  NAND2X1 U1708 ( .A(arr[813]), .B(n1221), .Y(n3202) );
  OAI21X1 U1709 ( .A(n2319), .B(n1220), .C(n3203), .Y(n4291) );
  NAND2X1 U1710 ( .A(arr[814]), .B(n1221), .Y(n3203) );
  OAI21X1 U1711 ( .A(n2321), .B(n1220), .C(n3204), .Y(n4292) );
  NAND2X1 U1712 ( .A(arr[815]), .B(n1221), .Y(n3204) );
  OAI21X1 U1714 ( .A(n1335), .B(n1218), .C(n3206), .Y(n4293) );
  NAND2X1 U1715 ( .A(arr[816]), .B(n1219), .Y(n3206) );
  OAI21X1 U1716 ( .A(n1334), .B(n1218), .C(n3207), .Y(n4294) );
  NAND2X1 U1717 ( .A(arr[817]), .B(n1219), .Y(n3207) );
  OAI21X1 U1718 ( .A(n1333), .B(n1218), .C(n3208), .Y(n4295) );
  NAND2X1 U1719 ( .A(arr[818]), .B(n1218), .Y(n3208) );
  OAI21X1 U1720 ( .A(n1332), .B(n1218), .C(n3209), .Y(n4296) );
  NAND2X1 U1721 ( .A(arr[819]), .B(n1218), .Y(n3209) );
  OAI21X1 U1722 ( .A(n1331), .B(n1218), .C(n3210), .Y(n4297) );
  NAND2X1 U1723 ( .A(arr[820]), .B(n1219), .Y(n3210) );
  OAI21X1 U1724 ( .A(n1330), .B(n1218), .C(n3211), .Y(n4298) );
  NAND2X1 U1725 ( .A(arr[821]), .B(n1219), .Y(n3211) );
  OAI21X1 U1726 ( .A(n1329), .B(n1218), .C(n3212), .Y(n4299) );
  NAND2X1 U1727 ( .A(arr[822]), .B(n1219), .Y(n3212) );
  OAI21X1 U1728 ( .A(n1328), .B(n1218), .C(n3213), .Y(n4300) );
  NAND2X1 U1729 ( .A(arr[823]), .B(n1219), .Y(n3213) );
  OAI21X1 U1730 ( .A(n1327), .B(n1218), .C(n3214), .Y(n4301) );
  NAND2X1 U1731 ( .A(arr[824]), .B(n1219), .Y(n3214) );
  OAI21X1 U1732 ( .A(n1326), .B(n1219), .C(n3215), .Y(n4302) );
  NAND2X1 U1733 ( .A(arr[825]), .B(n1219), .Y(n3215) );
  OAI21X1 U1734 ( .A(n1325), .B(n1219), .C(n3216), .Y(n4303) );
  NAND2X1 U1735 ( .A(arr[826]), .B(n1219), .Y(n3216) );
  OAI21X1 U1736 ( .A(n1324), .B(n1219), .C(n3217), .Y(n4304) );
  NAND2X1 U1737 ( .A(arr[827]), .B(n1219), .Y(n3217) );
  OAI21X1 U1738 ( .A(n1323), .B(n1218), .C(n3218), .Y(n4305) );
  NAND2X1 U1739 ( .A(arr[828]), .B(n1219), .Y(n3218) );
  OAI21X1 U1740 ( .A(n1322), .B(n1218), .C(n3219), .Y(n4306) );
  NAND2X1 U1741 ( .A(arr[829]), .B(n1219), .Y(n3219) );
  OAI21X1 U1742 ( .A(n1321), .B(n1218), .C(n3220), .Y(n4307) );
  NAND2X1 U1743 ( .A(arr[830]), .B(n1219), .Y(n3220) );
  OAI21X1 U1744 ( .A(n1320), .B(n1218), .C(n3221), .Y(n4308) );
  NAND2X1 U1745 ( .A(arr[831]), .B(n1219), .Y(n3221) );
  AND2X1 U1747 ( .A(n3187), .B(n2944), .Y(n2640) );
  OAI21X1 U1748 ( .A(n2291), .B(n1216), .C(n3223), .Y(n4309) );
  NAND2X1 U1749 ( .A(arr[832]), .B(n1217), .Y(n3223) );
  OAI21X1 U1750 ( .A(n2293), .B(n1216), .C(n3224), .Y(n4310) );
  NAND2X1 U1751 ( .A(arr[833]), .B(n1217), .Y(n3224) );
  OAI21X1 U1752 ( .A(n2295), .B(n1216), .C(n3225), .Y(n4311) );
  NAND2X1 U1753 ( .A(arr[834]), .B(n1216), .Y(n3225) );
  OAI21X1 U1754 ( .A(n2297), .B(n1216), .C(n3226), .Y(n4312) );
  NAND2X1 U1755 ( .A(arr[835]), .B(n1216), .Y(n3226) );
  OAI21X1 U1756 ( .A(n2299), .B(n1216), .C(n3227), .Y(n4313) );
  NAND2X1 U1757 ( .A(arr[836]), .B(n1217), .Y(n3227) );
  OAI21X1 U1758 ( .A(n2301), .B(n1216), .C(n3228), .Y(n4314) );
  NAND2X1 U1759 ( .A(arr[837]), .B(n1217), .Y(n3228) );
  OAI21X1 U1760 ( .A(n2303), .B(n1216), .C(n3229), .Y(n4315) );
  NAND2X1 U1761 ( .A(arr[838]), .B(n1217), .Y(n3229) );
  OAI21X1 U1762 ( .A(n2305), .B(n1216), .C(n3230), .Y(n4316) );
  NAND2X1 U1763 ( .A(arr[839]), .B(n1217), .Y(n3230) );
  OAI21X1 U1764 ( .A(n2307), .B(n1216), .C(n3231), .Y(n4317) );
  NAND2X1 U1765 ( .A(arr[840]), .B(n1217), .Y(n3231) );
  OAI21X1 U1766 ( .A(n2309), .B(n1217), .C(n3232), .Y(n4318) );
  NAND2X1 U1767 ( .A(arr[841]), .B(n1217), .Y(n3232) );
  OAI21X1 U1768 ( .A(n2311), .B(n1217), .C(n3233), .Y(n4319) );
  NAND2X1 U1769 ( .A(arr[842]), .B(n1217), .Y(n3233) );
  OAI21X1 U1770 ( .A(n2313), .B(n1217), .C(n3234), .Y(n4320) );
  NAND2X1 U1771 ( .A(arr[843]), .B(n1217), .Y(n3234) );
  OAI21X1 U1772 ( .A(n2315), .B(n1216), .C(n3235), .Y(n4321) );
  NAND2X1 U1773 ( .A(arr[844]), .B(n1217), .Y(n3235) );
  OAI21X1 U1774 ( .A(n2317), .B(n1216), .C(n3236), .Y(n4322) );
  NAND2X1 U1775 ( .A(arr[845]), .B(n1217), .Y(n3236) );
  OAI21X1 U1776 ( .A(n2319), .B(n1216), .C(n3237), .Y(n4323) );
  NAND2X1 U1777 ( .A(arr[846]), .B(n1217), .Y(n3237) );
  OAI21X1 U1778 ( .A(n2321), .B(n1216), .C(n3238), .Y(n4324) );
  NAND2X1 U1779 ( .A(arr[847]), .B(n1217), .Y(n3238) );
  OAI21X1 U1781 ( .A(n2291), .B(n1214), .C(n3240), .Y(n4325) );
  NAND2X1 U1782 ( .A(arr[848]), .B(n1215), .Y(n3240) );
  OAI21X1 U1783 ( .A(n2293), .B(n1214), .C(n3241), .Y(n4326) );
  NAND2X1 U1784 ( .A(arr[849]), .B(n1215), .Y(n3241) );
  OAI21X1 U1785 ( .A(n2295), .B(n1214), .C(n3242), .Y(n4327) );
  NAND2X1 U1786 ( .A(arr[850]), .B(n1214), .Y(n3242) );
  OAI21X1 U1787 ( .A(n2297), .B(n1214), .C(n3243), .Y(n4328) );
  NAND2X1 U1788 ( .A(arr[851]), .B(n1214), .Y(n3243) );
  OAI21X1 U1789 ( .A(n2299), .B(n1214), .C(n3244), .Y(n4329) );
  NAND2X1 U1790 ( .A(arr[852]), .B(n1215), .Y(n3244) );
  OAI21X1 U1791 ( .A(n2301), .B(n1214), .C(n3245), .Y(n4330) );
  NAND2X1 U1792 ( .A(arr[853]), .B(n1215), .Y(n3245) );
  OAI21X1 U1793 ( .A(n2303), .B(n1214), .C(n3246), .Y(n4331) );
  NAND2X1 U1794 ( .A(arr[854]), .B(n1215), .Y(n3246) );
  OAI21X1 U1795 ( .A(n2305), .B(n1214), .C(n3247), .Y(n4332) );
  NAND2X1 U1796 ( .A(arr[855]), .B(n1215), .Y(n3247) );
  OAI21X1 U1797 ( .A(n2307), .B(n1214), .C(n3248), .Y(n4333) );
  NAND2X1 U1798 ( .A(arr[856]), .B(n1215), .Y(n3248) );
  OAI21X1 U1799 ( .A(n2309), .B(n1215), .C(n3249), .Y(n4334) );
  NAND2X1 U1800 ( .A(arr[857]), .B(n1215), .Y(n3249) );
  OAI21X1 U1801 ( .A(n2311), .B(n1215), .C(n3250), .Y(n4335) );
  NAND2X1 U1802 ( .A(arr[858]), .B(n1215), .Y(n3250) );
  OAI21X1 U1803 ( .A(n2313), .B(n1215), .C(n3251), .Y(n4336) );
  NAND2X1 U1804 ( .A(arr[859]), .B(n1215), .Y(n3251) );
  OAI21X1 U1805 ( .A(n2315), .B(n1214), .C(n3252), .Y(n4337) );
  NAND2X1 U1806 ( .A(arr[860]), .B(n1215), .Y(n3252) );
  OAI21X1 U1807 ( .A(n2317), .B(n1214), .C(n3253), .Y(n4338) );
  NAND2X1 U1808 ( .A(arr[861]), .B(n1215), .Y(n3253) );
  OAI21X1 U1809 ( .A(n2319), .B(n1214), .C(n3254), .Y(n4339) );
  NAND2X1 U1810 ( .A(arr[862]), .B(n1215), .Y(n3254) );
  OAI21X1 U1811 ( .A(n2321), .B(n1214), .C(n3255), .Y(n4340) );
  NAND2X1 U1812 ( .A(arr[863]), .B(n1215), .Y(n3255) );
  AND2X1 U1814 ( .A(n3187), .B(n2979), .Y(n2675) );
  OAI21X1 U1815 ( .A(n2291), .B(n1212), .C(n3257), .Y(n4341) );
  NAND2X1 U1816 ( .A(arr[864]), .B(n1213), .Y(n3257) );
  OAI21X1 U1817 ( .A(n2293), .B(n1212), .C(n3258), .Y(n4342) );
  NAND2X1 U1818 ( .A(arr[865]), .B(n1213), .Y(n3258) );
  OAI21X1 U1819 ( .A(n2295), .B(n1212), .C(n3259), .Y(n4343) );
  NAND2X1 U1820 ( .A(arr[866]), .B(n1212), .Y(n3259) );
  OAI21X1 U1821 ( .A(n2297), .B(n1212), .C(n3260), .Y(n4344) );
  NAND2X1 U1822 ( .A(arr[867]), .B(n1212), .Y(n3260) );
  OAI21X1 U1823 ( .A(n2299), .B(n1212), .C(n3261), .Y(n4345) );
  NAND2X1 U1824 ( .A(arr[868]), .B(n1213), .Y(n3261) );
  OAI21X1 U1825 ( .A(n2301), .B(n1212), .C(n3262), .Y(n4346) );
  NAND2X1 U1826 ( .A(arr[869]), .B(n1213), .Y(n3262) );
  OAI21X1 U1827 ( .A(n2303), .B(n1212), .C(n3263), .Y(n4347) );
  NAND2X1 U1828 ( .A(arr[870]), .B(n1213), .Y(n3263) );
  OAI21X1 U1829 ( .A(n2305), .B(n1212), .C(n3264), .Y(n4348) );
  NAND2X1 U1830 ( .A(arr[871]), .B(n1213), .Y(n3264) );
  OAI21X1 U1831 ( .A(n2307), .B(n1212), .C(n3265), .Y(n4349) );
  NAND2X1 U1832 ( .A(arr[872]), .B(n1213), .Y(n3265) );
  OAI21X1 U1833 ( .A(n2309), .B(n1213), .C(n3266), .Y(n4350) );
  NAND2X1 U1834 ( .A(arr[873]), .B(n1213), .Y(n3266) );
  OAI21X1 U1835 ( .A(n2311), .B(n1213), .C(n3267), .Y(n4351) );
  NAND2X1 U1836 ( .A(arr[874]), .B(n1213), .Y(n3267) );
  OAI21X1 U1837 ( .A(n2313), .B(n1213), .C(n3268), .Y(n4352) );
  NAND2X1 U1838 ( .A(arr[875]), .B(n1213), .Y(n3268) );
  OAI21X1 U1839 ( .A(n2315), .B(n1212), .C(n3269), .Y(n4353) );
  NAND2X1 U1840 ( .A(arr[876]), .B(n1213), .Y(n3269) );
  OAI21X1 U1841 ( .A(n2317), .B(n1212), .C(n3270), .Y(n4354) );
  NAND2X1 U1842 ( .A(arr[877]), .B(n1213), .Y(n3270) );
  OAI21X1 U1843 ( .A(n2319), .B(n1212), .C(n3271), .Y(n4355) );
  NAND2X1 U1844 ( .A(arr[878]), .B(n1213), .Y(n3271) );
  OAI21X1 U1845 ( .A(n2321), .B(n1212), .C(n3272), .Y(n4356) );
  NAND2X1 U1846 ( .A(arr[879]), .B(n1213), .Y(n3272) );
  OAI21X1 U1848 ( .A(n2291), .B(n1210), .C(n3274), .Y(n4357) );
  NAND2X1 U1849 ( .A(arr[880]), .B(n1211), .Y(n3274) );
  OAI21X1 U1850 ( .A(n2293), .B(n1210), .C(n3275), .Y(n4358) );
  NAND2X1 U1851 ( .A(arr[881]), .B(n1211), .Y(n3275) );
  OAI21X1 U1852 ( .A(n2295), .B(n1210), .C(n3276), .Y(n4359) );
  NAND2X1 U1853 ( .A(arr[882]), .B(n1210), .Y(n3276) );
  OAI21X1 U1854 ( .A(n2297), .B(n1210), .C(n3277), .Y(n4360) );
  NAND2X1 U1855 ( .A(arr[883]), .B(n1210), .Y(n3277) );
  OAI21X1 U1856 ( .A(n2299), .B(n1210), .C(n3278), .Y(n4361) );
  NAND2X1 U1857 ( .A(arr[884]), .B(n1211), .Y(n3278) );
  OAI21X1 U1858 ( .A(n2301), .B(n1210), .C(n3279), .Y(n4362) );
  NAND2X1 U1859 ( .A(arr[885]), .B(n1211), .Y(n3279) );
  OAI21X1 U1860 ( .A(n2303), .B(n1210), .C(n3280), .Y(n4363) );
  NAND2X1 U1861 ( .A(arr[886]), .B(n1211), .Y(n3280) );
  OAI21X1 U1862 ( .A(n2305), .B(n1210), .C(n3281), .Y(n4364) );
  NAND2X1 U1863 ( .A(arr[887]), .B(n1211), .Y(n3281) );
  OAI21X1 U1864 ( .A(n2307), .B(n1210), .C(n3282), .Y(n4365) );
  NAND2X1 U1865 ( .A(arr[888]), .B(n1211), .Y(n3282) );
  OAI21X1 U1866 ( .A(n2309), .B(n1211), .C(n3283), .Y(n4366) );
  NAND2X1 U1867 ( .A(arr[889]), .B(n1211), .Y(n3283) );
  OAI21X1 U1868 ( .A(n2311), .B(n1211), .C(n3284), .Y(n4367) );
  NAND2X1 U1869 ( .A(arr[890]), .B(n1211), .Y(n3284) );
  OAI21X1 U1870 ( .A(n2313), .B(n1211), .C(n3285), .Y(n4368) );
  NAND2X1 U1871 ( .A(arr[891]), .B(n1211), .Y(n3285) );
  OAI21X1 U1872 ( .A(n2315), .B(n1210), .C(n3286), .Y(n4369) );
  NAND2X1 U1873 ( .A(arr[892]), .B(n1211), .Y(n3286) );
  OAI21X1 U1874 ( .A(n2317), .B(n1210), .C(n3287), .Y(n4370) );
  NAND2X1 U1875 ( .A(arr[893]), .B(n1211), .Y(n3287) );
  OAI21X1 U1876 ( .A(n2319), .B(n1210), .C(n3288), .Y(n4371) );
  NAND2X1 U1877 ( .A(arr[894]), .B(n1211), .Y(n3288) );
  OAI21X1 U1878 ( .A(n2321), .B(n1210), .C(n3289), .Y(n4372) );
  NAND2X1 U1879 ( .A(arr[895]), .B(n1211), .Y(n3289) );
  AND2X1 U1881 ( .A(n3187), .B(n3014), .Y(n2710) );
  NOR2X1 U1882 ( .A(n3290), .B(wr_ptr[3]), .Y(n3187) );
  OAI21X1 U1883 ( .A(n2291), .B(n1208), .C(n3292), .Y(n4373) );
  NAND2X1 U1884 ( .A(arr[896]), .B(n1209), .Y(n3292) );
  OAI21X1 U1885 ( .A(n2293), .B(n1208), .C(n3293), .Y(n4374) );
  NAND2X1 U1886 ( .A(arr[897]), .B(n1209), .Y(n3293) );
  OAI21X1 U1887 ( .A(n2295), .B(n1208), .C(n3294), .Y(n4375) );
  NAND2X1 U1888 ( .A(arr[898]), .B(n1208), .Y(n3294) );
  OAI21X1 U1889 ( .A(n2297), .B(n1208), .C(n3295), .Y(n4376) );
  NAND2X1 U1890 ( .A(arr[899]), .B(n1208), .Y(n3295) );
  OAI21X1 U1891 ( .A(n2299), .B(n1208), .C(n3296), .Y(n4377) );
  NAND2X1 U1892 ( .A(arr[900]), .B(n1209), .Y(n3296) );
  OAI21X1 U1893 ( .A(n2301), .B(n1208), .C(n3297), .Y(n4378) );
  NAND2X1 U1894 ( .A(arr[901]), .B(n1209), .Y(n3297) );
  OAI21X1 U1895 ( .A(n2303), .B(n1208), .C(n3298), .Y(n4379) );
  NAND2X1 U1896 ( .A(arr[902]), .B(n1209), .Y(n3298) );
  OAI21X1 U1897 ( .A(n2305), .B(n1208), .C(n3299), .Y(n4380) );
  NAND2X1 U1898 ( .A(arr[903]), .B(n1209), .Y(n3299) );
  OAI21X1 U1899 ( .A(n2307), .B(n1208), .C(n3300), .Y(n4381) );
  NAND2X1 U1900 ( .A(arr[904]), .B(n1209), .Y(n3300) );
  OAI21X1 U1901 ( .A(n2309), .B(n1209), .C(n3301), .Y(n4382) );
  NAND2X1 U1902 ( .A(arr[905]), .B(n1209), .Y(n3301) );
  OAI21X1 U1903 ( .A(n2311), .B(n1209), .C(n3302), .Y(n4383) );
  NAND2X1 U1904 ( .A(arr[906]), .B(n1209), .Y(n3302) );
  OAI21X1 U1905 ( .A(n2313), .B(n1209), .C(n3303), .Y(n4384) );
  NAND2X1 U1906 ( .A(arr[907]), .B(n1209), .Y(n3303) );
  OAI21X1 U1907 ( .A(n2315), .B(n1208), .C(n3304), .Y(n4385) );
  NAND2X1 U1908 ( .A(arr[908]), .B(n1209), .Y(n3304) );
  OAI21X1 U1909 ( .A(n2317), .B(n1208), .C(n3305), .Y(n4386) );
  NAND2X1 U1910 ( .A(arr[909]), .B(n1209), .Y(n3305) );
  OAI21X1 U1911 ( .A(n2319), .B(n1208), .C(n3306), .Y(n4387) );
  NAND2X1 U1912 ( .A(arr[910]), .B(n1209), .Y(n3306) );
  OAI21X1 U1913 ( .A(n2321), .B(n1208), .C(n3307), .Y(n4388) );
  NAND2X1 U1914 ( .A(arr[911]), .B(n1209), .Y(n3307) );
  OAI21X1 U1916 ( .A(n2291), .B(n1206), .C(n3309), .Y(n4389) );
  NAND2X1 U1917 ( .A(arr[912]), .B(n1207), .Y(n3309) );
  OAI21X1 U1918 ( .A(n2293), .B(n1206), .C(n3310), .Y(n4390) );
  NAND2X1 U1919 ( .A(arr[913]), .B(n1207), .Y(n3310) );
  OAI21X1 U1920 ( .A(n2295), .B(n1206), .C(n3311), .Y(n4391) );
  NAND2X1 U1921 ( .A(arr[914]), .B(n1206), .Y(n3311) );
  OAI21X1 U1922 ( .A(n2297), .B(n1206), .C(n3312), .Y(n4392) );
  NAND2X1 U1923 ( .A(arr[915]), .B(n1206), .Y(n3312) );
  OAI21X1 U1924 ( .A(n2299), .B(n1206), .C(n3313), .Y(n4393) );
  NAND2X1 U1925 ( .A(arr[916]), .B(n1207), .Y(n3313) );
  OAI21X1 U1926 ( .A(n2301), .B(n1206), .C(n3314), .Y(n4394) );
  NAND2X1 U1927 ( .A(arr[917]), .B(n1207), .Y(n3314) );
  OAI21X1 U1928 ( .A(n2303), .B(n1206), .C(n3315), .Y(n4395) );
  NAND2X1 U1929 ( .A(arr[918]), .B(n1207), .Y(n3315) );
  OAI21X1 U1930 ( .A(n2305), .B(n1206), .C(n3316), .Y(n4396) );
  NAND2X1 U1931 ( .A(arr[919]), .B(n1207), .Y(n3316) );
  OAI21X1 U1932 ( .A(n2307), .B(n1206), .C(n3317), .Y(n4397) );
  NAND2X1 U1933 ( .A(arr[920]), .B(n1207), .Y(n3317) );
  OAI21X1 U1934 ( .A(n2309), .B(n1207), .C(n3318), .Y(n4398) );
  NAND2X1 U1935 ( .A(arr[921]), .B(n1207), .Y(n3318) );
  OAI21X1 U1936 ( .A(n2311), .B(n1207), .C(n3319), .Y(n4399) );
  NAND2X1 U1937 ( .A(arr[922]), .B(n1207), .Y(n3319) );
  OAI21X1 U1938 ( .A(n2313), .B(n1207), .C(n3320), .Y(n4400) );
  NAND2X1 U1939 ( .A(arr[923]), .B(n1207), .Y(n3320) );
  OAI21X1 U1940 ( .A(n2315), .B(n1206), .C(n3321), .Y(n4401) );
  NAND2X1 U1941 ( .A(arr[924]), .B(n1207), .Y(n3321) );
  OAI21X1 U1942 ( .A(n2317), .B(n1206), .C(n3322), .Y(n4402) );
  NAND2X1 U1943 ( .A(arr[925]), .B(n1207), .Y(n3322) );
  OAI21X1 U1944 ( .A(n2319), .B(n1206), .C(n3323), .Y(n4403) );
  NAND2X1 U1945 ( .A(arr[926]), .B(n1207), .Y(n3323) );
  OAI21X1 U1946 ( .A(n2321), .B(n1206), .C(n3324), .Y(n4404) );
  NAND2X1 U1947 ( .A(arr[927]), .B(n1207), .Y(n3324) );
  AND2X1 U1949 ( .A(n3325), .B(n2909), .Y(n2745) );
  NOR2X1 U1950 ( .A(wr_ptr[1]), .B(wr_ptr[2]), .Y(n2909) );
  OAI21X1 U1951 ( .A(n1335), .B(n1204), .C(n3327), .Y(n4405) );
  NAND2X1 U1952 ( .A(arr[928]), .B(n1205), .Y(n3327) );
  OAI21X1 U1953 ( .A(n1334), .B(n1204), .C(n3328), .Y(n4406) );
  NAND2X1 U1954 ( .A(arr[929]), .B(n1205), .Y(n3328) );
  OAI21X1 U1955 ( .A(n1333), .B(n1204), .C(n3329), .Y(n4407) );
  NAND2X1 U1956 ( .A(arr[930]), .B(n1204), .Y(n3329) );
  OAI21X1 U1957 ( .A(n1332), .B(n1204), .C(n3330), .Y(n4408) );
  NAND2X1 U1958 ( .A(arr[931]), .B(n1204), .Y(n3330) );
  OAI21X1 U1959 ( .A(n1331), .B(n1204), .C(n3331), .Y(n4409) );
  NAND2X1 U1960 ( .A(arr[932]), .B(n1205), .Y(n3331) );
  OAI21X1 U1961 ( .A(n1330), .B(n1204), .C(n3332), .Y(n4410) );
  NAND2X1 U1962 ( .A(arr[933]), .B(n1205), .Y(n3332) );
  OAI21X1 U1963 ( .A(n1329), .B(n1204), .C(n3333), .Y(n4411) );
  NAND2X1 U1964 ( .A(arr[934]), .B(n1205), .Y(n3333) );
  OAI21X1 U1965 ( .A(n1328), .B(n1204), .C(n3334), .Y(n4412) );
  NAND2X1 U1966 ( .A(arr[935]), .B(n1205), .Y(n3334) );
  OAI21X1 U1967 ( .A(n1327), .B(n1204), .C(n3335), .Y(n4413) );
  NAND2X1 U1968 ( .A(arr[936]), .B(n1205), .Y(n3335) );
  OAI21X1 U1969 ( .A(n1326), .B(n1205), .C(n3336), .Y(n4414) );
  NAND2X1 U1970 ( .A(arr[937]), .B(n1205), .Y(n3336) );
  OAI21X1 U1971 ( .A(n1325), .B(n1205), .C(n3337), .Y(n4415) );
  NAND2X1 U1972 ( .A(arr[938]), .B(n1205), .Y(n3337) );
  OAI21X1 U1973 ( .A(n1324), .B(n1205), .C(n3338), .Y(n4416) );
  NAND2X1 U1974 ( .A(arr[939]), .B(n1205), .Y(n3338) );
  OAI21X1 U1975 ( .A(n1323), .B(n1204), .C(n3339), .Y(n4417) );
  NAND2X1 U1976 ( .A(arr[940]), .B(n1205), .Y(n3339) );
  OAI21X1 U1977 ( .A(n1322), .B(n1204), .C(n3340), .Y(n4418) );
  NAND2X1 U1978 ( .A(arr[941]), .B(n1205), .Y(n3340) );
  OAI21X1 U1979 ( .A(n1321), .B(n1204), .C(n3341), .Y(n4419) );
  NAND2X1 U1980 ( .A(arr[942]), .B(n1205), .Y(n3341) );
  OAI21X1 U1981 ( .A(n1320), .B(n1204), .C(n3342), .Y(n4420) );
  NAND2X1 U1982 ( .A(arr[943]), .B(n1205), .Y(n3342) );
  OAI21X1 U1984 ( .A(n2291), .B(n1202), .C(n3344), .Y(n4421) );
  NAND2X1 U1985 ( .A(arr[944]), .B(n1203), .Y(n3344) );
  OAI21X1 U1986 ( .A(n2293), .B(n1202), .C(n3345), .Y(n4422) );
  NAND2X1 U1987 ( .A(arr[945]), .B(n1203), .Y(n3345) );
  OAI21X1 U1988 ( .A(n2295), .B(n1202), .C(n3346), .Y(n4423) );
  NAND2X1 U1989 ( .A(arr[946]), .B(n1202), .Y(n3346) );
  OAI21X1 U1990 ( .A(n2297), .B(n1202), .C(n3347), .Y(n4424) );
  NAND2X1 U1991 ( .A(arr[947]), .B(n1202), .Y(n3347) );
  OAI21X1 U1992 ( .A(n2299), .B(n1202), .C(n3348), .Y(n4425) );
  NAND2X1 U1993 ( .A(arr[948]), .B(n1203), .Y(n3348) );
  OAI21X1 U1994 ( .A(n2301), .B(n1202), .C(n3349), .Y(n4426) );
  NAND2X1 U1995 ( .A(arr[949]), .B(n1203), .Y(n3349) );
  OAI21X1 U1996 ( .A(n2303), .B(n1202), .C(n3350), .Y(n4427) );
  NAND2X1 U1997 ( .A(arr[950]), .B(n1203), .Y(n3350) );
  OAI21X1 U1998 ( .A(n2305), .B(n1202), .C(n3351), .Y(n4428) );
  NAND2X1 U1999 ( .A(arr[951]), .B(n1203), .Y(n3351) );
  OAI21X1 U2000 ( .A(n2307), .B(n1202), .C(n3352), .Y(n4429) );
  NAND2X1 U2001 ( .A(arr[952]), .B(n1203), .Y(n3352) );
  OAI21X1 U2002 ( .A(n2309), .B(n1203), .C(n3353), .Y(n4430) );
  NAND2X1 U2003 ( .A(arr[953]), .B(n1203), .Y(n3353) );
  OAI21X1 U2004 ( .A(n2311), .B(n1203), .C(n3354), .Y(n4431) );
  NAND2X1 U2005 ( .A(arr[954]), .B(n1203), .Y(n3354) );
  OAI21X1 U2006 ( .A(n2313), .B(n1203), .C(n3355), .Y(n4432) );
  NAND2X1 U2007 ( .A(arr[955]), .B(n1203), .Y(n3355) );
  OAI21X1 U2008 ( .A(n2315), .B(n1202), .C(n3356), .Y(n4433) );
  NAND2X1 U2009 ( .A(arr[956]), .B(n1203), .Y(n3356) );
  OAI21X1 U2010 ( .A(n2317), .B(n1202), .C(n3357), .Y(n4434) );
  NAND2X1 U2011 ( .A(arr[957]), .B(n1203), .Y(n3357) );
  OAI21X1 U2012 ( .A(n2319), .B(n1202), .C(n3358), .Y(n4435) );
  NAND2X1 U2013 ( .A(arr[958]), .B(n1203), .Y(n3358) );
  OAI21X1 U2014 ( .A(n2321), .B(n1202), .C(n3359), .Y(n4436) );
  NAND2X1 U2015 ( .A(arr[959]), .B(n1203), .Y(n3359) );
  AND2X1 U2017 ( .A(n3325), .B(n2944), .Y(n2780) );
  NOR2X1 U2018 ( .A(n3360), .B(wr_ptr[2]), .Y(n2944) );
  OAI21X1 U2019 ( .A(n1335), .B(n1200), .C(n3362), .Y(n4437) );
  NAND2X1 U2020 ( .A(arr[960]), .B(n1201), .Y(n3362) );
  OAI21X1 U2021 ( .A(n1334), .B(n1200), .C(n3363), .Y(n4438) );
  NAND2X1 U2022 ( .A(arr[961]), .B(n1201), .Y(n3363) );
  OAI21X1 U2023 ( .A(n1333), .B(n1200), .C(n3364), .Y(n4439) );
  NAND2X1 U2024 ( .A(arr[962]), .B(n1200), .Y(n3364) );
  OAI21X1 U2025 ( .A(n1332), .B(n1200), .C(n3365), .Y(n4440) );
  NAND2X1 U2026 ( .A(arr[963]), .B(n1200), .Y(n3365) );
  OAI21X1 U2027 ( .A(n1331), .B(n1200), .C(n3366), .Y(n4441) );
  NAND2X1 U2028 ( .A(arr[964]), .B(n1201), .Y(n3366) );
  OAI21X1 U2029 ( .A(n1330), .B(n1200), .C(n3367), .Y(n4442) );
  NAND2X1 U2030 ( .A(arr[965]), .B(n1201), .Y(n3367) );
  OAI21X1 U2031 ( .A(n1329), .B(n1200), .C(n3368), .Y(n4443) );
  NAND2X1 U2032 ( .A(arr[966]), .B(n1201), .Y(n3368) );
  OAI21X1 U2033 ( .A(n1328), .B(n1200), .C(n3369), .Y(n4444) );
  NAND2X1 U2034 ( .A(arr[967]), .B(n1201), .Y(n3369) );
  OAI21X1 U2035 ( .A(n1327), .B(n1200), .C(n3370), .Y(n4445) );
  NAND2X1 U2036 ( .A(arr[968]), .B(n1201), .Y(n3370) );
  OAI21X1 U2037 ( .A(n1326), .B(n1201), .C(n3371), .Y(n4446) );
  NAND2X1 U2038 ( .A(arr[969]), .B(n1201), .Y(n3371) );
  OAI21X1 U2039 ( .A(n1325), .B(n1201), .C(n3372), .Y(n4447) );
  NAND2X1 U2040 ( .A(arr[970]), .B(n1201), .Y(n3372) );
  OAI21X1 U2041 ( .A(n1324), .B(n1201), .C(n3373), .Y(n4448) );
  NAND2X1 U2042 ( .A(arr[971]), .B(n1201), .Y(n3373) );
  OAI21X1 U2043 ( .A(n1323), .B(n1200), .C(n3374), .Y(n4449) );
  NAND2X1 U2044 ( .A(arr[972]), .B(n1201), .Y(n3374) );
  OAI21X1 U2045 ( .A(n1322), .B(n1200), .C(n3375), .Y(n4450) );
  NAND2X1 U2046 ( .A(arr[973]), .B(n1201), .Y(n3375) );
  OAI21X1 U2047 ( .A(n1321), .B(n1200), .C(n3376), .Y(n4451) );
  NAND2X1 U2048 ( .A(arr[974]), .B(n1201), .Y(n3376) );
  OAI21X1 U2049 ( .A(n1320), .B(n1200), .C(n3377), .Y(n4452) );
  NAND2X1 U2050 ( .A(arr[975]), .B(n1201), .Y(n3377) );
  OAI21X1 U2052 ( .A(n2291), .B(n1198), .C(n3379), .Y(n4453) );
  NAND2X1 U2053 ( .A(arr[976]), .B(n1199), .Y(n3379) );
  OAI21X1 U2054 ( .A(n2293), .B(n1198), .C(n3380), .Y(n4454) );
  NAND2X1 U2055 ( .A(arr[977]), .B(n1199), .Y(n3380) );
  OAI21X1 U2056 ( .A(n2295), .B(n1198), .C(n3381), .Y(n4455) );
  NAND2X1 U2057 ( .A(arr[978]), .B(n1198), .Y(n3381) );
  OAI21X1 U2058 ( .A(n2297), .B(n1198), .C(n3382), .Y(n4456) );
  NAND2X1 U2059 ( .A(arr[979]), .B(n1198), .Y(n3382) );
  OAI21X1 U2060 ( .A(n2299), .B(n1198), .C(n3383), .Y(n4457) );
  NAND2X1 U2061 ( .A(arr[980]), .B(n1199), .Y(n3383) );
  OAI21X1 U2062 ( .A(n2301), .B(n1198), .C(n3384), .Y(n4458) );
  NAND2X1 U2063 ( .A(arr[981]), .B(n1199), .Y(n3384) );
  OAI21X1 U2064 ( .A(n2303), .B(n1198), .C(n3385), .Y(n4459) );
  NAND2X1 U2065 ( .A(arr[982]), .B(n1199), .Y(n3385) );
  OAI21X1 U2066 ( .A(n2305), .B(n1198), .C(n3386), .Y(n4460) );
  NAND2X1 U2067 ( .A(arr[983]), .B(n1199), .Y(n3386) );
  OAI21X1 U2068 ( .A(n2307), .B(n1198), .C(n3387), .Y(n4461) );
  NAND2X1 U2069 ( .A(arr[984]), .B(n1199), .Y(n3387) );
  OAI21X1 U2070 ( .A(n2309), .B(n1199), .C(n3388), .Y(n4462) );
  NAND2X1 U2071 ( .A(arr[985]), .B(n1199), .Y(n3388) );
  OAI21X1 U2072 ( .A(n2311), .B(n1199), .C(n3389), .Y(n4463) );
  NAND2X1 U2073 ( .A(arr[986]), .B(n1199), .Y(n3389) );
  OAI21X1 U2074 ( .A(n2313), .B(n1199), .C(n3390), .Y(n4464) );
  NAND2X1 U2075 ( .A(arr[987]), .B(n1199), .Y(n3390) );
  OAI21X1 U2076 ( .A(n2315), .B(n1198), .C(n3391), .Y(n4465) );
  NAND2X1 U2077 ( .A(arr[988]), .B(n1199), .Y(n3391) );
  OAI21X1 U2078 ( .A(n2317), .B(n1198), .C(n3392), .Y(n4466) );
  NAND2X1 U2079 ( .A(arr[989]), .B(n1199), .Y(n3392) );
  OAI21X1 U2080 ( .A(n2319), .B(n1198), .C(n3393), .Y(n4467) );
  NAND2X1 U2081 ( .A(arr[990]), .B(n1199), .Y(n3393) );
  OAI21X1 U2082 ( .A(n2321), .B(n1198), .C(n3394), .Y(n4468) );
  NAND2X1 U2083 ( .A(arr[991]), .B(n1199), .Y(n3394) );
  AND2X1 U2085 ( .A(n3325), .B(n2979), .Y(n2815) );
  NOR2X1 U2086 ( .A(n3395), .B(wr_ptr[1]), .Y(n2979) );
  OAI21X1 U2087 ( .A(n1335), .B(n1196), .C(n3397), .Y(n4469) );
  NAND2X1 U2088 ( .A(arr[992]), .B(n1197), .Y(n3397) );
  OAI21X1 U2089 ( .A(n1334), .B(n1196), .C(n3398), .Y(n4470) );
  NAND2X1 U2090 ( .A(arr[993]), .B(n1197), .Y(n3398) );
  OAI21X1 U2091 ( .A(n1333), .B(n1196), .C(n3399), .Y(n4471) );
  NAND2X1 U2092 ( .A(arr[994]), .B(n1196), .Y(n3399) );
  OAI21X1 U2093 ( .A(n1332), .B(n1196), .C(n3400), .Y(n4472) );
  NAND2X1 U2094 ( .A(arr[995]), .B(n1196), .Y(n3400) );
  OAI21X1 U2095 ( .A(n1331), .B(n1196), .C(n3401), .Y(n4473) );
  NAND2X1 U2096 ( .A(arr[996]), .B(n1197), .Y(n3401) );
  OAI21X1 U2097 ( .A(n1330), .B(n1196), .C(n3402), .Y(n4474) );
  NAND2X1 U2098 ( .A(arr[997]), .B(n1197), .Y(n3402) );
  OAI21X1 U2099 ( .A(n1329), .B(n1196), .C(n3403), .Y(n4475) );
  NAND2X1 U2100 ( .A(arr[998]), .B(n1197), .Y(n3403) );
  OAI21X1 U2101 ( .A(n1328), .B(n1196), .C(n3404), .Y(n4476) );
  NAND2X1 U2102 ( .A(arr[999]), .B(n1197), .Y(n3404) );
  OAI21X1 U2103 ( .A(n1327), .B(n1196), .C(n3405), .Y(n4477) );
  NAND2X1 U2104 ( .A(arr[1000]), .B(n1197), .Y(n3405) );
  OAI21X1 U2105 ( .A(n1326), .B(n1197), .C(n3406), .Y(n4478) );
  NAND2X1 U2106 ( .A(arr[1001]), .B(n1197), .Y(n3406) );
  OAI21X1 U2107 ( .A(n1325), .B(n1197), .C(n3407), .Y(n4479) );
  NAND2X1 U2108 ( .A(arr[1002]), .B(n1197), .Y(n3407) );
  OAI21X1 U2109 ( .A(n1324), .B(n1197), .C(n3408), .Y(n4480) );
  NAND2X1 U2110 ( .A(arr[1003]), .B(n1197), .Y(n3408) );
  OAI21X1 U2111 ( .A(n1323), .B(n1196), .C(n3409), .Y(n4481) );
  NAND2X1 U2112 ( .A(arr[1004]), .B(n1197), .Y(n3409) );
  OAI21X1 U2113 ( .A(n1322), .B(n1196), .C(n3410), .Y(n4482) );
  NAND2X1 U2114 ( .A(arr[1005]), .B(n1197), .Y(n3410) );
  OAI21X1 U2115 ( .A(n1321), .B(n1196), .C(n3411), .Y(n4483) );
  NAND2X1 U2116 ( .A(arr[1006]), .B(n1197), .Y(n3411) );
  OAI21X1 U2117 ( .A(n1320), .B(n1196), .C(n3412), .Y(n4484) );
  NAND2X1 U2118 ( .A(arr[1007]), .B(n1197), .Y(n3412) );
  OAI21X1 U2121 ( .A(n2291), .B(n1194), .C(n3415), .Y(n4485) );
  NAND2X1 U2122 ( .A(arr[1008]), .B(n1195), .Y(n3415) );
  OAI21X1 U2124 ( .A(n2293), .B(n1194), .C(n3416), .Y(n4486) );
  NAND2X1 U2125 ( .A(arr[1009]), .B(n1195), .Y(n3416) );
  OAI21X1 U2127 ( .A(n2295), .B(n1194), .C(n3417), .Y(n4487) );
  NAND2X1 U2128 ( .A(arr[1010]), .B(n1194), .Y(n3417) );
  OAI21X1 U2130 ( .A(n2297), .B(n1194), .C(n3418), .Y(n4488) );
  NAND2X1 U2131 ( .A(arr[1011]), .B(n1194), .Y(n3418) );
  OAI21X1 U2133 ( .A(n2299), .B(n1194), .C(n3419), .Y(n4489) );
  NAND2X1 U2134 ( .A(arr[1012]), .B(n1195), .Y(n3419) );
  OAI21X1 U2136 ( .A(n2301), .B(n1194), .C(n3420), .Y(n4490) );
  NAND2X1 U2137 ( .A(arr[1013]), .B(n1195), .Y(n3420) );
  OAI21X1 U2139 ( .A(n2303), .B(n1194), .C(n3421), .Y(n4491) );
  NAND2X1 U2140 ( .A(arr[1014]), .B(n1195), .Y(n3421) );
  OAI21X1 U2142 ( .A(n2305), .B(n1194), .C(n3422), .Y(n4492) );
  NAND2X1 U2143 ( .A(arr[1015]), .B(n1195), .Y(n3422) );
  OAI21X1 U2145 ( .A(n2307), .B(n1194), .C(n3423), .Y(n4493) );
  NAND2X1 U2146 ( .A(arr[1016]), .B(n1195), .Y(n3423) );
  OAI21X1 U2148 ( .A(n2309), .B(n1195), .C(n3424), .Y(n4494) );
  NAND2X1 U2149 ( .A(arr[1017]), .B(n1195), .Y(n3424) );
  OAI21X1 U2151 ( .A(n2311), .B(n1195), .C(n3425), .Y(n4495) );
  NAND2X1 U2152 ( .A(arr[1018]), .B(n1195), .Y(n3425) );
  OAI21X1 U2154 ( .A(n2313), .B(n1195), .C(n3426), .Y(n4496) );
  NAND2X1 U2155 ( .A(arr[1019]), .B(n1195), .Y(n3426) );
  OAI21X1 U2157 ( .A(n2315), .B(n1194), .C(n3427), .Y(n4497) );
  NAND2X1 U2158 ( .A(arr[1020]), .B(n1195), .Y(n3427) );
  OAI21X1 U2160 ( .A(n2317), .B(n1194), .C(n3428), .Y(n4498) );
  NAND2X1 U2161 ( .A(arr[1021]), .B(n1195), .Y(n3428) );
  OAI21X1 U2163 ( .A(n2319), .B(n1194), .C(n3429), .Y(n4499) );
  NAND2X1 U2164 ( .A(arr[1022]), .B(n1195), .Y(n3429) );
  OAI21X1 U2166 ( .A(n2321), .B(n1194), .C(n3430), .Y(n4500) );
  NAND2X1 U2167 ( .A(arr[1023]), .B(n1195), .Y(n3430) );
  AND2X1 U2169 ( .A(n3325), .B(n3014), .Y(n2850) );
  NOR2X1 U2170 ( .A(n3395), .B(n3360), .Y(n3014) );
  NOR2X1 U2171 ( .A(n3290), .B(n3152), .Y(n3325) );
  AND2X1 U2173 ( .A(wr_ptr[5]), .B(n2870), .Y(n3413) );
  OAI21X1 U2175 ( .A(n2871), .B(n3431), .C(n3432), .Y(n4501) );
  NAND2X1 U2176 ( .A(n91), .B(n2870), .Y(n3432) );
  OAI21X1 U2178 ( .A(n3290), .B(n3431), .C(n3433), .Y(n4502) );
  NAND2X1 U2179 ( .A(n90), .B(n2870), .Y(n3433) );
  OAI21X1 U2181 ( .A(n3152), .B(n3431), .C(n3434), .Y(n4503) );
  NAND2X1 U2182 ( .A(n89), .B(n2870), .Y(n3434) );
  OAI21X1 U2184 ( .A(n3395), .B(n3431), .C(n3435), .Y(n4504) );
  NAND2X1 U2185 ( .A(n88), .B(n2870), .Y(n3435) );
  OAI21X1 U2187 ( .A(n3360), .B(n3431), .C(n3436), .Y(n4505) );
  NAND2X1 U2188 ( .A(n87), .B(n2870), .Y(n3436) );
  OAI21X1 U2190 ( .A(n2852), .B(n3431), .C(n3437), .Y(n4506) );
  NAND2X1 U2191 ( .A(n86), .B(n2870), .Y(n3437) );
  NAND2X1 U2193 ( .A(n3438), .B(n3439), .Y(n3431) );
  OAI21X1 U2196 ( .A(n3441), .B(n3442), .C(n3443), .Y(n4507) );
  AOI22X1 U2197 ( .A(n97), .B(n3444), .C(n1136), .D(n3445), .Y(n3443) );
  OAI21X1 U2199 ( .A(n3441), .B(n3446), .C(n3447), .Y(n4508) );
  AOI22X1 U2200 ( .A(n96), .B(n3444), .C(n1135), .D(n3445), .Y(n3447) );
  OAI21X1 U2201 ( .A(n3441), .B(n3448), .C(n3449), .Y(n4509) );
  AOI22X1 U2202 ( .A(n95), .B(n3444), .C(n1134), .D(n3445), .Y(n3449) );
  OAI21X1 U2203 ( .A(n3441), .B(n3450), .C(n3451), .Y(n4510) );
  AOI22X1 U2204 ( .A(n94), .B(n3444), .C(n1133), .D(n3445), .Y(n3451) );
  OAI21X1 U2205 ( .A(n3441), .B(n3452), .C(n3453), .Y(n4511) );
  AOI22X1 U2206 ( .A(n98), .B(n3444), .C(n1137), .D(n3445), .Y(n3453) );
  OAI21X1 U2208 ( .A(n3441), .B(n3454), .C(n3455), .Y(n4512) );
  AOI22X1 U2209 ( .A(n93), .B(n3444), .C(n1132), .D(n3445), .Y(n3455) );
  OAI21X1 U2210 ( .A(n3441), .B(n3456), .C(n3457), .Y(n4513) );
  AOI22X1 U2211 ( .A(n92), .B(n3444), .C(n1131), .D(n3445), .Y(n3457) );
  NAND3X1 U2213 ( .A(n3441), .B(get), .C(n3459), .Y(n3458) );
  NOR2X1 U2214 ( .A(reset), .B(empty), .Y(n3459) );
  NOR2X1 U2215 ( .A(n3460), .B(n2289), .Y(n3444) );
  OAI21X1 U2217 ( .A(n3440), .B(n2289), .C(n3461), .Y(n3460) );
  NAND3X1 U2218 ( .A(n3462), .B(n3439), .C(n3463), .Y(n3461) );
  NOR2X1 U2219 ( .A(n3464), .B(n3465), .Y(n3463) );
  AOI21X1 U2221 ( .A(n3467), .B(n3468), .C(n3469), .Y(n3466) );
  OAI21X1 U2222 ( .A(empty), .B(n3464), .C(n3439), .Y(n2289) );
  NOR2X1 U2225 ( .A(n3465), .B(full), .Y(n3440) );
  NOR2X1 U2227 ( .A(n3468), .B(n3469), .Y(full) );
  NAND3X1 U2228 ( .A(fillcount[1]), .B(n3456), .C(fillcount[2]), .Y(n3468) );
  NOR2X1 U2229 ( .A(n3469), .B(n3467), .Y(empty) );
  NAND3X1 U2230 ( .A(n3454), .B(n3450), .C(n3456), .Y(n3467) );
  NAND3X1 U2234 ( .A(n3448), .B(n3446), .C(n3470), .Y(n3469) );
  NOR2X1 U2235 ( .A(fillcount[6]), .B(fillcount[5]), .Y(n3470) );
  INVX2 U3 ( .A(n2281), .Y(n3471) );
  INVX2 U5 ( .A(n2284), .Y(n3472) );
  INVX2 U7 ( .A(n2285), .Y(n3473) );
  INVX2 U9 ( .A(n2286), .Y(n3474) );
  INVX2 U11 ( .A(n2287), .Y(n3475) );
  INVX2 U13 ( .A(n2288), .Y(n3476) );
  INVX2 U16 ( .A(n2289), .Y(n2283) );
  INVX2 U2123 ( .A(data_in[0]), .Y(n2291) );
  INVX2 U2126 ( .A(data_in[1]), .Y(n2293) );
  INVX2 U2129 ( .A(data_in[2]), .Y(n2295) );
  INVX2 U2132 ( .A(data_in[3]), .Y(n2297) );
  INVX2 U2135 ( .A(data_in[4]), .Y(n2299) );
  INVX2 U2138 ( .A(data_in[5]), .Y(n2301) );
  INVX2 U2141 ( .A(data_in[6]), .Y(n2303) );
  INVX2 U2144 ( .A(data_in[7]), .Y(n2305) );
  INVX2 U2147 ( .A(data_in[8]), .Y(n2307) );
  INVX2 U2150 ( .A(data_in[9]), .Y(n2309) );
  INVX2 U2153 ( .A(data_in[10]), .Y(n2311) );
  INVX2 U2156 ( .A(data_in[11]), .Y(n2313) );
  INVX2 U2159 ( .A(data_in[12]), .Y(n2315) );
  INVX2 U2162 ( .A(data_in[13]), .Y(n2317) );
  INVX2 U2165 ( .A(data_in[14]), .Y(n2319) );
  INVX2 U2174 ( .A(data_in[15]), .Y(n2321) );
  INVX2 U2177 ( .A(wr_ptr[5]), .Y(n2871) );
  INVX2 U2180 ( .A(wr_ptr[4]), .Y(n3290) );
  INVX2 U2183 ( .A(wr_ptr[3]), .Y(n3152) );
  INVX2 U2186 ( .A(wr_ptr[2]), .Y(n3395) );
  INVX2 U2189 ( .A(wr_ptr[1]), .Y(n3360) );
  INVX2 U2195 ( .A(wr_ptr[0]), .Y(n2852) );
  INVX2 U2207 ( .A(fillcount[6]), .Y(n3452) );
  INVX2 U2212 ( .A(n3458), .Y(n3445) );
  INVX2 U2216 ( .A(n3460), .Y(n3441) );
  INVX2 U2220 ( .A(n3466), .Y(n3462) );
  INVX2 U2223 ( .A(reset), .Y(n3439) );
  INVX2 U2224 ( .A(get), .Y(n3464) );
  INVX2 U2226 ( .A(put), .Y(n3465) );
  INVX2 U2232 ( .A(fillcount[2]), .Y(n3450) );
  INVX2 U2233 ( .A(fillcount[1]), .Y(n3454) );
  INVX2 U2236 ( .A(fillcount[4]), .Y(n3446) );
  INVX2 U2237 ( .A(fillcount[3]), .Y(n3448) );
  FIFO_DEPTH_P26_WIDTH16_DW01_dec_0 sub_55 ( .A(fillcount), .SUM({n1137, n1136, 
        n1135, n1134, n1133, n1132, n1131}) );
  FIFO_DEPTH_P26_WIDTH16_DW01_inc_0 add_54 ( .A({n18, n17, n16, n15, n14, n13}), .SUM({n1130, n1129, n1128, n1127, n1126, n1125}) );
  FIFO_DEPTH_P26_WIDTH16_DW01_inc_1 add_50 ( .A(fillcount), .SUM({n98, n97, 
        n96, n95, n94, n93, n92}) );
  FIFO_DEPTH_P26_WIDTH16_DW01_inc_2 add_49 ( .A(wr_ptr), .SUM({n91, n90, n89, 
        n88, n87, n86}) );
  AND2X2 U49 ( .A(n2850), .B(n2342), .Y(n1) );
  AND2X2 U82 ( .A(n2815), .B(n2342), .Y(n2) );
  AND2X2 U115 ( .A(n2780), .B(n2342), .Y(n3) );
  AND2X2 U148 ( .A(n2745), .B(n2342), .Y(n4) );
  AND2X2 U181 ( .A(n2710), .B(n2342), .Y(n5) );
  AND2X2 U214 ( .A(n2675), .B(n2342), .Y(n6) );
  AND2X2 U247 ( .A(n2640), .B(n2342), .Y(n7) );
  AND2X2 U280 ( .A(n2605), .B(n2342), .Y(n8) );
  AND2X2 U313 ( .A(n2570), .B(n2342), .Y(n9) );
  AND2X2 U346 ( .A(n2535), .B(n2342), .Y(n10) );
  AND2X2 U379 ( .A(n2500), .B(n2342), .Y(n11) );
  AND2X2 U412 ( .A(n2465), .B(n2342), .Y(n12) );
  AND2X2 U445 ( .A(n2430), .B(n2342), .Y(n19) );
  AND2X2 U478 ( .A(n2395), .B(n2342), .Y(n20) );
  AND2X2 U511 ( .A(n2360), .B(n2342), .Y(n21) );
  AND2X2 U544 ( .A(n2850), .B(n2323), .Y(n22) );
  AND2X2 U577 ( .A(n2815), .B(n2323), .Y(n23) );
  AND2X2 U610 ( .A(n2780), .B(n2323), .Y(n24) );
  AND2X2 U643 ( .A(n2745), .B(n2323), .Y(n25) );
  AND2X2 U676 ( .A(n2710), .B(n2323), .Y(n26) );
  AND2X2 U709 ( .A(n2675), .B(n2323), .Y(n27) );
  AND2X2 U742 ( .A(n2640), .B(n2323), .Y(n28) );
  AND2X2 U775 ( .A(n2605), .B(n2323), .Y(n29) );
  AND2X2 U808 ( .A(n2570), .B(n2323), .Y(n30) );
  AND2X2 U841 ( .A(n2535), .B(n2323), .Y(n31) );
  AND2X2 U874 ( .A(n2500), .B(n2323), .Y(n32) );
  AND2X2 U907 ( .A(n2465), .B(n2323), .Y(n33) );
  AND2X2 U940 ( .A(n2430), .B(n2323), .Y(n34) );
  AND2X2 U973 ( .A(n2395), .B(n2323), .Y(n35) );
  AND2X2 U1006 ( .A(n2360), .B(n2323), .Y(n36) );
  AND2X2 U1039 ( .A(n2342), .B(n2324), .Y(n37) );
  AND2X2 U1040 ( .A(n2323), .B(n2324), .Y(n38) );
  AND2X2 U1073 ( .A(n2907), .B(n2850), .Y(n39) );
  AND2X2 U1074 ( .A(n2907), .B(n2815), .Y(n40) );
  AND2X2 U1108 ( .A(n2907), .B(n2780), .Y(n41) );
  AND2X2 U1141 ( .A(n2907), .B(n2745), .Y(n42) );
  AND2X2 U1175 ( .A(n2907), .B(n2710), .Y(n43) );
  AND2X2 U1208 ( .A(n2907), .B(n2675), .Y(n44) );
  AND2X2 U1242 ( .A(n2907), .B(n2640), .Y(n45) );
  AND2X2 U1275 ( .A(n2907), .B(n2605), .Y(n46) );
  AND2X2 U1309 ( .A(n2907), .B(n2570), .Y(n47) );
  AND2X2 U1342 ( .A(n2907), .B(n2535), .Y(n48) );
  AND2X2 U1377 ( .A(n2907), .B(n2500), .Y(n49) );
  AND2X2 U1410 ( .A(n2907), .B(n2465), .Y(n50) );
  AND2X2 U1444 ( .A(n2907), .B(n2430), .Y(n51) );
  AND2X2 U1477 ( .A(n2907), .B(n2395), .Y(n52) );
  AND2X2 U1511 ( .A(n2907), .B(n2360), .Y(n53) );
  AND2X2 U1544 ( .A(n2907), .B(n2324), .Y(n54) );
  AND2X2 U1578 ( .A(n2889), .B(n2850), .Y(n55) );
  AND2X2 U1611 ( .A(n2889), .B(n2815), .Y(n56) );
  AND2X2 U1646 ( .A(n2889), .B(n2780), .Y(n57) );
  AND2X2 U1679 ( .A(n2889), .B(n2745), .Y(n58) );
  AND2X2 U1713 ( .A(n2889), .B(n2710), .Y(n59) );
  AND2X2 U1746 ( .A(n2889), .B(n2675), .Y(n60) );
  AND2X2 U1780 ( .A(n2889), .B(n2640), .Y(n61) );
  AND2X2 U1813 ( .A(n2889), .B(n2605), .Y(n62) );
  AND2X2 U1847 ( .A(n2889), .B(n2570), .Y(n63) );
  AND2X2 U1880 ( .A(n2889), .B(n2535), .Y(n64) );
  AND2X2 U1915 ( .A(n2889), .B(n2500), .Y(n65) );
  AND2X2 U1948 ( .A(n2889), .B(n2465), .Y(n66) );
  AND2X2 U1983 ( .A(n2889), .B(n2430), .Y(n67) );
  AND2X2 U2016 ( .A(n2889), .B(n2395), .Y(n68) );
  AND2X2 U2051 ( .A(n2889), .B(n2360), .Y(n69) );
  AND2X2 U2084 ( .A(n2889), .B(n2324), .Y(n70) );
  INVX2 U2119 ( .A(n70), .Y(n1256) );
  INVX2 U2120 ( .A(n69), .Y(n1252) );
  INVX2 U2168 ( .A(n68), .Y(n1248) );
  INVX2 U2172 ( .A(n67), .Y(n1244) );
  INVX2 U2192 ( .A(n66), .Y(n1240) );
  INVX2 U2194 ( .A(n65), .Y(n1236) );
  INVX2 U2198 ( .A(n64), .Y(n1232) );
  INVX2 U2231 ( .A(n63), .Y(n1228) );
  INVX2 U2238 ( .A(n62), .Y(n1224) );
  INVX2 U2239 ( .A(n61), .Y(n1220) );
  INVX2 U2240 ( .A(n60), .Y(n1216) );
  INVX2 U2241 ( .A(n59), .Y(n1212) );
  INVX2 U2242 ( .A(n58), .Y(n1208) );
  INVX2 U2243 ( .A(n57), .Y(n1204) );
  INVX2 U2244 ( .A(n56), .Y(n1200) );
  INVX2 U2245 ( .A(n55), .Y(n1196) );
  INVX2 U2246 ( .A(n70), .Y(n1257) );
  INVX2 U2247 ( .A(n69), .Y(n1253) );
  INVX2 U2248 ( .A(n68), .Y(n1249) );
  INVX2 U2249 ( .A(n67), .Y(n1245) );
  INVX2 U2250 ( .A(n66), .Y(n1241) );
  INVX2 U2251 ( .A(n65), .Y(n1237) );
  INVX2 U2252 ( .A(n64), .Y(n1233) );
  INVX2 U2253 ( .A(n63), .Y(n1229) );
  INVX2 U2254 ( .A(n62), .Y(n1225) );
  INVX2 U2255 ( .A(n61), .Y(n1221) );
  INVX2 U2256 ( .A(n60), .Y(n1217) );
  INVX2 U2257 ( .A(n59), .Y(n1213) );
  INVX2 U2258 ( .A(n58), .Y(n1209) );
  INVX2 U2259 ( .A(n57), .Y(n1205) );
  INVX2 U2260 ( .A(n56), .Y(n1201) );
  INVX2 U2261 ( .A(n55), .Y(n1197) );
  INVX2 U2262 ( .A(n36), .Y(n1317) );
  INVX2 U2263 ( .A(n35), .Y(n1313) );
  INVX2 U2264 ( .A(n34), .Y(n1309) );
  INVX2 U2265 ( .A(n33), .Y(n1305) );
  INVX2 U2266 ( .A(n32), .Y(n1301) );
  INVX2 U2267 ( .A(n31), .Y(n1297) );
  INVX2 U2268 ( .A(n30), .Y(n1293) );
  INVX2 U2269 ( .A(n29), .Y(n1289) );
  INVX2 U2270 ( .A(n28), .Y(n1285) );
  INVX2 U2271 ( .A(n27), .Y(n1281) );
  INVX2 U2272 ( .A(n26), .Y(n1277) );
  INVX2 U2273 ( .A(n25), .Y(n1273) );
  INVX2 U2274 ( .A(n24), .Y(n1269) );
  INVX2 U2275 ( .A(n23), .Y(n1265) );
  INVX2 U2276 ( .A(n22), .Y(n1261) );
  INVX2 U2277 ( .A(n38), .Y(n1337) );
  INVX2 U2278 ( .A(n37), .Y(n1318) );
  INVX2 U2279 ( .A(n54), .Y(n1254) );
  INVX2 U2280 ( .A(n53), .Y(n1250) );
  INVX2 U2281 ( .A(n52), .Y(n1246) );
  INVX2 U2282 ( .A(n51), .Y(n1242) );
  INVX2 U2283 ( .A(n50), .Y(n1238) );
  INVX2 U2284 ( .A(n49), .Y(n1234) );
  INVX2 U2285 ( .A(n48), .Y(n1230) );
  INVX2 U2286 ( .A(n47), .Y(n1226) );
  INVX2 U2287 ( .A(n46), .Y(n1222) );
  INVX2 U2288 ( .A(n45), .Y(n1218) );
  INVX2 U2289 ( .A(n44), .Y(n1214) );
  INVX2 U2290 ( .A(n43), .Y(n1210) );
  INVX2 U2291 ( .A(n42), .Y(n1206) );
  INVX2 U2292 ( .A(n41), .Y(n1202) );
  INVX2 U2293 ( .A(n40), .Y(n1198) );
  INVX2 U2294 ( .A(n39), .Y(n1194) );
  INVX2 U2295 ( .A(n37), .Y(n1319) );
  INVX2 U2296 ( .A(n54), .Y(n1255) );
  INVX2 U2297 ( .A(n53), .Y(n1251) );
  INVX2 U2298 ( .A(n52), .Y(n1247) );
  INVX2 U2299 ( .A(n51), .Y(n1243) );
  INVX2 U2300 ( .A(n50), .Y(n1239) );
  INVX2 U2301 ( .A(n49), .Y(n1235) );
  INVX2 U2302 ( .A(n48), .Y(n1231) );
  INVX2 U2303 ( .A(n47), .Y(n1227) );
  INVX2 U2304 ( .A(n46), .Y(n1223) );
  INVX2 U2305 ( .A(n45), .Y(n1219) );
  INVX2 U2306 ( .A(n44), .Y(n1215) );
  INVX2 U2307 ( .A(n43), .Y(n1211) );
  INVX2 U2308 ( .A(n42), .Y(n1207) );
  INVX2 U2309 ( .A(n41), .Y(n1203) );
  INVX2 U2310 ( .A(n40), .Y(n1199) );
  INVX2 U2311 ( .A(n39), .Y(n1195) );
  INVX2 U2312 ( .A(n21), .Y(n1315) );
  INVX2 U2313 ( .A(n20), .Y(n1311) );
  INVX2 U2314 ( .A(n19), .Y(n1307) );
  INVX2 U2315 ( .A(n12), .Y(n1303) );
  INVX2 U2316 ( .A(n11), .Y(n1299) );
  INVX2 U2317 ( .A(n10), .Y(n1295) );
  INVX2 U2318 ( .A(n9), .Y(n1291) );
  INVX2 U2319 ( .A(n8), .Y(n1287) );
  INVX2 U2320 ( .A(n7), .Y(n1283) );
  INVX2 U2321 ( .A(n6), .Y(n1279) );
  INVX2 U2322 ( .A(n5), .Y(n1275) );
  INVX2 U2323 ( .A(n4), .Y(n1271) );
  INVX2 U2324 ( .A(n3), .Y(n1267) );
  INVX2 U2325 ( .A(n2), .Y(n1263) );
  INVX2 U2326 ( .A(n1), .Y(n1259) );
  INVX2 U2327 ( .A(n36), .Y(n1316) );
  INVX2 U2328 ( .A(n35), .Y(n1312) );
  INVX2 U2329 ( .A(n34), .Y(n1308) );
  INVX2 U2330 ( .A(n33), .Y(n1304) );
  INVX2 U2331 ( .A(n32), .Y(n1300) );
  INVX2 U2332 ( .A(n31), .Y(n1296) );
  INVX2 U2333 ( .A(n30), .Y(n1292) );
  INVX2 U2334 ( .A(n29), .Y(n1288) );
  INVX2 U2335 ( .A(n28), .Y(n1284) );
  INVX2 U2336 ( .A(n27), .Y(n1280) );
  INVX2 U2337 ( .A(n26), .Y(n1276) );
  INVX2 U2338 ( .A(n25), .Y(n1272) );
  INVX2 U2339 ( .A(n24), .Y(n1268) );
  INVX2 U2340 ( .A(n23), .Y(n1264) );
  INVX2 U2341 ( .A(n22), .Y(n1260) );
  INVX2 U2342 ( .A(n38), .Y(n1336) );
  INVX2 U2343 ( .A(n21), .Y(n1314) );
  INVX2 U2344 ( .A(n20), .Y(n1310) );
  INVX2 U2345 ( .A(n19), .Y(n1306) );
  INVX2 U2346 ( .A(n12), .Y(n1302) );
  INVX2 U2347 ( .A(n11), .Y(n1298) );
  INVX2 U2348 ( .A(n10), .Y(n1294) );
  INVX2 U2349 ( .A(n9), .Y(n1290) );
  INVX2 U2350 ( .A(n8), .Y(n1286) );
  INVX2 U2351 ( .A(n7), .Y(n1282) );
  INVX2 U2352 ( .A(n6), .Y(n1278) );
  INVX2 U2353 ( .A(n5), .Y(n1274) );
  INVX2 U2354 ( .A(n4), .Y(n1270) );
  INVX2 U2355 ( .A(n3), .Y(n1266) );
  INVX2 U2356 ( .A(n2), .Y(n1262) );
  INVX2 U2357 ( .A(n1), .Y(n1258) );
  INVX2 U2358 ( .A(data_in[0]), .Y(n1335) );
  INVX2 U2359 ( .A(data_in[1]), .Y(n1334) );
  INVX2 U2360 ( .A(data_in[2]), .Y(n1333) );
  INVX2 U2361 ( .A(data_in[3]), .Y(n1332) );
  INVX2 U2362 ( .A(data_in[4]), .Y(n1331) );
  INVX2 U2363 ( .A(data_in[5]), .Y(n1330) );
  INVX2 U2364 ( .A(data_in[6]), .Y(n1329) );
  INVX2 U2365 ( .A(data_in[7]), .Y(n1328) );
  INVX2 U2366 ( .A(data_in[8]), .Y(n1327) );
  INVX2 U2367 ( .A(data_in[9]), .Y(n1326) );
  INVX2 U2368 ( .A(data_in[10]), .Y(n1325) );
  INVX2 U2369 ( .A(data_in[11]), .Y(n1324) );
  INVX2 U2370 ( .A(data_in[12]), .Y(n1323) );
  INVX2 U2371 ( .A(data_in[13]), .Y(n1322) );
  INVX2 U2372 ( .A(data_in[14]), .Y(n1321) );
  INVX2 U2373 ( .A(data_in[15]), .Y(n1320) );
  BUFX2 U2374 ( .A(n1120), .Y(n1078) );
  BUFX2 U2375 ( .A(n1120), .Y(n1077) );
  BUFX2 U2376 ( .A(n1120), .Y(n1079) );
  BUFX2 U2377 ( .A(n1121), .Y(n1080) );
  BUFX2 U2378 ( .A(n1121), .Y(n1082) );
  BUFX2 U2379 ( .A(n1121), .Y(n1081) );
  BUFX2 U2380 ( .A(n1122), .Y(n1083) );
  BUFX2 U2381 ( .A(n1122), .Y(n1084) );
  BUFX2 U2382 ( .A(n1123), .Y(n1086) );
  BUFX2 U2383 ( .A(n1122), .Y(n1085) );
  BUFX2 U2384 ( .A(n1123), .Y(n1087) );
  BUFX2 U2385 ( .A(n1123), .Y(n1088) );
  BUFX2 U2386 ( .A(n1124), .Y(n1090) );
  BUFX2 U2387 ( .A(n1124), .Y(n1089) );
  BUFX2 U2388 ( .A(n1124), .Y(n1091) );
  BUFX2 U2389 ( .A(n1138), .Y(n1092) );
  BUFX2 U2390 ( .A(n1138), .Y(n1094) );
  BUFX2 U2391 ( .A(n1138), .Y(n1093) );
  BUFX2 U2392 ( .A(n1139), .Y(n1095) );
  BUFX2 U2393 ( .A(n1139), .Y(n1096) );
  BUFX2 U2394 ( .A(n1140), .Y(n1098) );
  BUFX2 U2395 ( .A(n1139), .Y(n1097) );
  BUFX2 U2396 ( .A(n1140), .Y(n1099) );
  BUFX2 U2397 ( .A(n1140), .Y(n1100) );
  BUFX2 U2398 ( .A(n1141), .Y(n1102) );
  BUFX2 U2399 ( .A(n1141), .Y(n1101) );
  BUFX2 U2400 ( .A(n1141), .Y(n1103) );
  BUFX2 U2401 ( .A(n1142), .Y(n1104) );
  BUFX2 U2402 ( .A(n1142), .Y(n1106) );
  BUFX2 U2403 ( .A(n1142), .Y(n1105) );
  BUFX2 U2404 ( .A(n1143), .Y(n1107) );
  BUFX2 U2405 ( .A(n1143), .Y(n1108) );
  BUFX2 U2406 ( .A(n1144), .Y(n1110) );
  BUFX2 U2407 ( .A(n1143), .Y(n1109) );
  BUFX2 U2408 ( .A(n1144), .Y(n1111) );
  BUFX2 U2409 ( .A(n1144), .Y(n1112) );
  BUFX2 U2410 ( .A(n1145), .Y(n1114) );
  BUFX2 U2411 ( .A(n1145), .Y(n1113) );
  BUFX2 U2412 ( .A(n1145), .Y(n1115) );
  BUFX2 U2413 ( .A(n1146), .Y(n1116) );
  BUFX2 U2414 ( .A(n1146), .Y(n1118) );
  BUFX2 U2415 ( .A(n1146), .Y(n1117) );
  BUFX2 U2416 ( .A(n1170), .Y(n1148) );
  BUFX2 U2417 ( .A(n1170), .Y(n1149) );
  BUFX2 U2418 ( .A(n1170), .Y(n1150) );
  BUFX2 U2419 ( .A(n1171), .Y(n1151) );
  BUFX2 U2420 ( .A(n1171), .Y(n1152) );
  BUFX2 U2421 ( .A(n1171), .Y(n1153) );
  BUFX2 U2422 ( .A(n1172), .Y(n1154) );
  BUFX2 U2423 ( .A(n1172), .Y(n1155) );
  BUFX2 U2424 ( .A(n1172), .Y(n1156) );
  BUFX2 U2425 ( .A(n1173), .Y(n1157) );
  BUFX2 U2426 ( .A(n1173), .Y(n1158) );
  BUFX2 U2427 ( .A(n1173), .Y(n1159) );
  BUFX2 U2428 ( .A(n1174), .Y(n1160) );
  BUFX2 U2429 ( .A(n1174), .Y(n1161) );
  BUFX2 U2430 ( .A(n1174), .Y(n1162) );
  BUFX2 U2431 ( .A(n1175), .Y(n1163) );
  BUFX2 U2432 ( .A(n1175), .Y(n1164) );
  BUFX2 U2433 ( .A(n1175), .Y(n1165) );
  BUFX2 U2434 ( .A(n1176), .Y(n1166) );
  BUFX2 U2435 ( .A(n1176), .Y(n1167) );
  BUFX2 U2436 ( .A(n1176), .Y(n1168) );
  BUFX2 U2437 ( .A(n15), .Y(n1178) );
  BUFX2 U2438 ( .A(n15), .Y(n1179) );
  BUFX2 U2439 ( .A(n15), .Y(n1180) );
  BUFX2 U2440 ( .A(n15), .Y(n1181) );
  BUFX2 U2441 ( .A(n15), .Y(n1182) );
  BUFX2 U2442 ( .A(n15), .Y(n1183) );
  BUFX2 U2443 ( .A(n15), .Y(n1184) );
  BUFX2 U2444 ( .A(n15), .Y(n1185) );
  BUFX2 U2445 ( .A(n15), .Y(n1186) );
  BUFX2 U2446 ( .A(n15), .Y(n1187) );
  BUFX2 U2447 ( .A(n15), .Y(n1177) );
  BUFX2 U2448 ( .A(n1119), .Y(n1076) );
  BUFX2 U2449 ( .A(n13), .Y(n1119) );
  BUFX2 U2450 ( .A(n13), .Y(n1120) );
  BUFX2 U2451 ( .A(n13), .Y(n1121) );
  BUFX2 U2452 ( .A(n13), .Y(n1122) );
  BUFX2 U2453 ( .A(n13), .Y(n1123) );
  BUFX2 U2454 ( .A(n13), .Y(n1124) );
  BUFX2 U2455 ( .A(n13), .Y(n1138) );
  BUFX2 U2456 ( .A(n13), .Y(n1139) );
  BUFX2 U2457 ( .A(n13), .Y(n1140) );
  BUFX2 U2458 ( .A(n13), .Y(n1141) );
  BUFX2 U2459 ( .A(n13), .Y(n1142) );
  BUFX2 U2460 ( .A(n13), .Y(n1143) );
  BUFX2 U2461 ( .A(n13), .Y(n1144) );
  BUFX2 U2462 ( .A(n13), .Y(n1145) );
  BUFX2 U2463 ( .A(n13), .Y(n1146) );
  INVX2 U2464 ( .A(fillcount[0]), .Y(n3456) );
  BUFX2 U2465 ( .A(n16), .Y(n1189) );
  BUFX2 U2466 ( .A(n16), .Y(n1190) );
  BUFX2 U2467 ( .A(n16), .Y(n1191) );
  BUFX2 U2468 ( .A(n16), .Y(n1192) );
  BUFX2 U2469 ( .A(n16), .Y(n1193) );
  BUFX2 U2470 ( .A(n16), .Y(n1188) );
  BUFX2 U2471 ( .A(n1169), .Y(n1147) );
  BUFX2 U2472 ( .A(n14), .Y(n1169) );
  BUFX2 U2473 ( .A(n14), .Y(n1170) );
  BUFX2 U2474 ( .A(n14), .Y(n1171) );
  BUFX2 U2475 ( .A(n14), .Y(n1172) );
  BUFX2 U2476 ( .A(n14), .Y(n1173) );
  BUFX2 U2477 ( .A(n14), .Y(n1174) );
  BUFX2 U2478 ( .A(n14), .Y(n1175) );
  BUFX2 U2479 ( .A(n14), .Y(n1176) );
  MUX2X1 U2480 ( .B(n72), .A(n73), .S(n1147), .Y(n71) );
  MUX2X1 U2481 ( .B(n75), .A(n76), .S(n1147), .Y(n74) );
  MUX2X1 U2482 ( .B(n78), .A(n79), .S(n1147), .Y(n77) );
  MUX2X1 U2483 ( .B(n81), .A(n82), .S(n1147), .Y(n80) );
  MUX2X1 U2484 ( .B(n84), .A(n85), .S(n1188), .Y(n83) );
  MUX2X1 U2485 ( .B(n100), .A(n101), .S(n1148), .Y(n99) );
  MUX2X1 U2486 ( .B(n103), .A(n104), .S(n1148), .Y(n102) );
  MUX2X1 U2487 ( .B(n106), .A(n107), .S(n1148), .Y(n105) );
  MUX2X1 U2488 ( .B(n109), .A(n110), .S(n1148), .Y(n108) );
  MUX2X1 U2489 ( .B(n112), .A(n113), .S(n1188), .Y(n111) );
  MUX2X1 U2490 ( .B(n115), .A(n116), .S(n1148), .Y(n114) );
  MUX2X1 U2491 ( .B(n118), .A(n119), .S(n1148), .Y(n117) );
  MUX2X1 U2492 ( .B(n121), .A(n122), .S(n1148), .Y(n120) );
  MUX2X1 U2493 ( .B(n124), .A(n125), .S(n1148), .Y(n123) );
  MUX2X1 U2494 ( .B(n127), .A(n128), .S(n1188), .Y(n126) );
  MUX2X1 U2495 ( .B(n130), .A(n131), .S(n1148), .Y(n129) );
  MUX2X1 U2496 ( .B(n133), .A(n134), .S(n1148), .Y(n132) );
  MUX2X1 U2497 ( .B(n136), .A(n137), .S(n1148), .Y(n135) );
  MUX2X1 U2498 ( .B(n139), .A(n140), .S(n1148), .Y(n138) );
  MUX2X1 U2499 ( .B(n142), .A(n143), .S(n1188), .Y(n141) );
  MUX2X1 U2500 ( .B(n144), .A(n145), .S(n18), .Y(data_out[0]) );
  MUX2X1 U2501 ( .B(n147), .A(n148), .S(n1149), .Y(n146) );
  MUX2X1 U2502 ( .B(n150), .A(n151), .S(n1149), .Y(n149) );
  MUX2X1 U2503 ( .B(n153), .A(n154), .S(n1149), .Y(n152) );
  MUX2X1 U2504 ( .B(n156), .A(n157), .S(n1149), .Y(n155) );
  MUX2X1 U2505 ( .B(n159), .A(n160), .S(n1189), .Y(n158) );
  MUX2X1 U2506 ( .B(n162), .A(n163), .S(n1149), .Y(n161) );
  MUX2X1 U2507 ( .B(n165), .A(n166), .S(n1149), .Y(n164) );
  MUX2X1 U2508 ( .B(n168), .A(n169), .S(n1149), .Y(n167) );
  MUX2X1 U2509 ( .B(n171), .A(n172), .S(n1149), .Y(n170) );
  MUX2X1 U2510 ( .B(n174), .A(n175), .S(n1189), .Y(n173) );
  MUX2X1 U2511 ( .B(n177), .A(n178), .S(n1149), .Y(n176) );
  MUX2X1 U2512 ( .B(n180), .A(n181), .S(n1149), .Y(n179) );
  MUX2X1 U2513 ( .B(n183), .A(n184), .S(n1149), .Y(n182) );
  MUX2X1 U2514 ( .B(n186), .A(n187), .S(n1149), .Y(n185) );
  MUX2X1 U2515 ( .B(n189), .A(n190), .S(n1189), .Y(n188) );
  MUX2X1 U2516 ( .B(n192), .A(n193), .S(n1150), .Y(n191) );
  MUX2X1 U2517 ( .B(n195), .A(n196), .S(n1150), .Y(n194) );
  MUX2X1 U2518 ( .B(n198), .A(n199), .S(n1150), .Y(n197) );
  MUX2X1 U2519 ( .B(n201), .A(n202), .S(n1150), .Y(n200) );
  MUX2X1 U2520 ( .B(n204), .A(n205), .S(n1189), .Y(n203) );
  MUX2X1 U2521 ( .B(n206), .A(n207), .S(n18), .Y(data_out[1]) );
  MUX2X1 U2522 ( .B(n209), .A(n210), .S(n1150), .Y(n208) );
  MUX2X1 U2523 ( .B(n212), .A(n213), .S(n1150), .Y(n211) );
  MUX2X1 U2524 ( .B(n215), .A(n216), .S(n1150), .Y(n214) );
  MUX2X1 U2525 ( .B(n218), .A(n219), .S(n1150), .Y(n217) );
  MUX2X1 U2526 ( .B(n221), .A(n222), .S(n1189), .Y(n220) );
  MUX2X1 U2527 ( .B(n224), .A(n225), .S(n1150), .Y(n223) );
  MUX2X1 U2528 ( .B(n227), .A(n228), .S(n1150), .Y(n226) );
  MUX2X1 U2529 ( .B(n230), .A(n231), .S(n1150), .Y(n229) );
  MUX2X1 U2530 ( .B(n233), .A(n234), .S(n1150), .Y(n232) );
  MUX2X1 U2531 ( .B(n236), .A(n237), .S(n1189), .Y(n235) );
  MUX2X1 U2532 ( .B(n239), .A(n240), .S(n1151), .Y(n238) );
  MUX2X1 U2533 ( .B(n242), .A(n243), .S(n1151), .Y(n241) );
  MUX2X1 U2534 ( .B(n245), .A(n246), .S(n1151), .Y(n244) );
  MUX2X1 U2535 ( .B(n248), .A(n249), .S(n1151), .Y(n247) );
  MUX2X1 U2536 ( .B(n251), .A(n252), .S(n1189), .Y(n250) );
  MUX2X1 U2537 ( .B(n254), .A(n255), .S(n1151), .Y(n253) );
  MUX2X1 U2538 ( .B(n257), .A(n258), .S(n1151), .Y(n256) );
  MUX2X1 U2539 ( .B(n260), .A(n261), .S(n1151), .Y(n259) );
  MUX2X1 U2540 ( .B(n263), .A(n264), .S(n1151), .Y(n262) );
  MUX2X1 U2541 ( .B(n266), .A(n267), .S(n1189), .Y(n265) );
  MUX2X1 U2542 ( .B(n268), .A(n269), .S(n18), .Y(data_out[2]) );
  MUX2X1 U2543 ( .B(n271), .A(n272), .S(n1151), .Y(n270) );
  MUX2X1 U2544 ( .B(n274), .A(n275), .S(n1151), .Y(n273) );
  MUX2X1 U2545 ( .B(n277), .A(n278), .S(n1151), .Y(n276) );
  MUX2X1 U2546 ( .B(n280), .A(n281), .S(n1151), .Y(n279) );
  MUX2X1 U2547 ( .B(n283), .A(n284), .S(n1189), .Y(n282) );
  MUX2X1 U2548 ( .B(n286), .A(n287), .S(n1152), .Y(n285) );
  MUX2X1 U2549 ( .B(n289), .A(n290), .S(n1152), .Y(n288) );
  MUX2X1 U2550 ( .B(n292), .A(n293), .S(n1152), .Y(n291) );
  MUX2X1 U2551 ( .B(n295), .A(n296), .S(n1152), .Y(n294) );
  MUX2X1 U2552 ( .B(n298), .A(n299), .S(n1189), .Y(n297) );
  MUX2X1 U2553 ( .B(n301), .A(n302), .S(n1152), .Y(n300) );
  MUX2X1 U2554 ( .B(n304), .A(n305), .S(n1152), .Y(n303) );
  MUX2X1 U2555 ( .B(n307), .A(n308), .S(n1152), .Y(n306) );
  MUX2X1 U2556 ( .B(n310), .A(n311), .S(n1152), .Y(n309) );
  MUX2X1 U2557 ( .B(n313), .A(n314), .S(n1189), .Y(n312) );
  MUX2X1 U2558 ( .B(n316), .A(n317), .S(n1152), .Y(n315) );
  MUX2X1 U2559 ( .B(n319), .A(n320), .S(n1152), .Y(n318) );
  MUX2X1 U2560 ( .B(n322), .A(n323), .S(n1152), .Y(n321) );
  MUX2X1 U2561 ( .B(n325), .A(n326), .S(n1152), .Y(n324) );
  MUX2X1 U2562 ( .B(n328), .A(n329), .S(n1189), .Y(n327) );
  MUX2X1 U2563 ( .B(n330), .A(n331), .S(n18), .Y(data_out[3]) );
  MUX2X1 U2564 ( .B(n333), .A(n334), .S(n1153), .Y(n332) );
  MUX2X1 U2565 ( .B(n336), .A(n337), .S(n1153), .Y(n335) );
  MUX2X1 U2566 ( .B(n339), .A(n340), .S(n1153), .Y(n338) );
  MUX2X1 U2567 ( .B(n342), .A(n343), .S(n1153), .Y(n341) );
  MUX2X1 U2568 ( .B(n345), .A(n346), .S(n1190), .Y(n344) );
  MUX2X1 U2569 ( .B(n348), .A(n349), .S(n1153), .Y(n347) );
  MUX2X1 U2570 ( .B(n351), .A(n352), .S(n1153), .Y(n350) );
  MUX2X1 U2571 ( .B(n354), .A(n355), .S(n1153), .Y(n353) );
  MUX2X1 U2572 ( .B(n357), .A(n358), .S(n1153), .Y(n356) );
  MUX2X1 U2573 ( .B(n360), .A(n361), .S(n1190), .Y(n359) );
  MUX2X1 U2574 ( .B(n363), .A(n364), .S(n1153), .Y(n362) );
  MUX2X1 U2575 ( .B(n366), .A(n367), .S(n1153), .Y(n365) );
  MUX2X1 U2576 ( .B(n369), .A(n370), .S(n1153), .Y(n368) );
  MUX2X1 U2577 ( .B(n372), .A(n373), .S(n1153), .Y(n371) );
  MUX2X1 U2578 ( .B(n375), .A(n376), .S(n1190), .Y(n374) );
  MUX2X1 U2579 ( .B(n378), .A(n379), .S(n1154), .Y(n377) );
  MUX2X1 U2580 ( .B(n381), .A(n382), .S(n1154), .Y(n380) );
  MUX2X1 U2581 ( .B(n384), .A(n385), .S(n1154), .Y(n383) );
  MUX2X1 U2582 ( .B(n387), .A(n388), .S(n1154), .Y(n386) );
  MUX2X1 U2583 ( .B(n390), .A(n391), .S(n1190), .Y(n389) );
  MUX2X1 U2584 ( .B(n392), .A(n393), .S(n18), .Y(data_out[4]) );
  MUX2X1 U2585 ( .B(n395), .A(n396), .S(n1154), .Y(n394) );
  MUX2X1 U2586 ( .B(n398), .A(n399), .S(n1154), .Y(n397) );
  MUX2X1 U2587 ( .B(n401), .A(n402), .S(n1154), .Y(n400) );
  MUX2X1 U2588 ( .B(n404), .A(n405), .S(n1154), .Y(n403) );
  MUX2X1 U2589 ( .B(n407), .A(n408), .S(n1190), .Y(n406) );
  MUX2X1 U2590 ( .B(n410), .A(n411), .S(n1154), .Y(n409) );
  MUX2X1 U2591 ( .B(n413), .A(n414), .S(n1154), .Y(n412) );
  MUX2X1 U2592 ( .B(n416), .A(n417), .S(n1154), .Y(n415) );
  MUX2X1 U2593 ( .B(n419), .A(n420), .S(n1154), .Y(n418) );
  MUX2X1 U2594 ( .B(n422), .A(n423), .S(n1190), .Y(n421) );
  MUX2X1 U2595 ( .B(n425), .A(n426), .S(n1155), .Y(n424) );
  MUX2X1 U2596 ( .B(n428), .A(n429), .S(n1155), .Y(n427) );
  MUX2X1 U2597 ( .B(n431), .A(n432), .S(n1155), .Y(n430) );
  MUX2X1 U2598 ( .B(n434), .A(n435), .S(n1155), .Y(n433) );
  MUX2X1 U2599 ( .B(n437), .A(n438), .S(n1190), .Y(n436) );
  MUX2X1 U2600 ( .B(n440), .A(n441), .S(n1155), .Y(n439) );
  MUX2X1 U2601 ( .B(n443), .A(n444), .S(n1155), .Y(n442) );
  MUX2X1 U2602 ( .B(n446), .A(n447), .S(n1155), .Y(n445) );
  MUX2X1 U2603 ( .B(n449), .A(n450), .S(n1155), .Y(n448) );
  MUX2X1 U2604 ( .B(n452), .A(n453), .S(n1190), .Y(n451) );
  MUX2X1 U2605 ( .B(n454), .A(n455), .S(n18), .Y(data_out[5]) );
  MUX2X1 U2606 ( .B(n457), .A(n458), .S(n1155), .Y(n456) );
  MUX2X1 U2607 ( .B(n460), .A(n461), .S(n1155), .Y(n459) );
  MUX2X1 U2608 ( .B(n463), .A(n464), .S(n1155), .Y(n462) );
  MUX2X1 U2609 ( .B(n466), .A(n467), .S(n1155), .Y(n465) );
  MUX2X1 U2610 ( .B(n469), .A(n470), .S(n1190), .Y(n468) );
  MUX2X1 U2611 ( .B(n472), .A(n473), .S(n1156), .Y(n471) );
  MUX2X1 U2612 ( .B(n475), .A(n476), .S(n1156), .Y(n474) );
  MUX2X1 U2613 ( .B(n478), .A(n479), .S(n1156), .Y(n477) );
  MUX2X1 U2614 ( .B(n481), .A(n482), .S(n1156), .Y(n480) );
  MUX2X1 U2615 ( .B(n484), .A(n485), .S(n1190), .Y(n483) );
  MUX2X1 U2616 ( .B(n487), .A(n488), .S(n1156), .Y(n486) );
  MUX2X1 U2617 ( .B(n490), .A(n491), .S(n1156), .Y(n489) );
  MUX2X1 U2618 ( .B(n493), .A(n494), .S(n1156), .Y(n492) );
  MUX2X1 U2619 ( .B(n496), .A(n497), .S(n1156), .Y(n495) );
  MUX2X1 U2620 ( .B(n499), .A(n500), .S(n1190), .Y(n498) );
  MUX2X1 U2621 ( .B(n502), .A(n503), .S(n1156), .Y(n501) );
  MUX2X1 U2622 ( .B(n505), .A(n506), .S(n1156), .Y(n504) );
  MUX2X1 U2623 ( .B(n508), .A(n509), .S(n1156), .Y(n507) );
  MUX2X1 U2624 ( .B(n511), .A(n512), .S(n1156), .Y(n510) );
  MUX2X1 U2625 ( .B(n514), .A(n515), .S(n1190), .Y(n513) );
  MUX2X1 U2626 ( .B(n516), .A(n517), .S(n18), .Y(data_out[6]) );
  MUX2X1 U2627 ( .B(n519), .A(n520), .S(n1157), .Y(n518) );
  MUX2X1 U2628 ( .B(n522), .A(n523), .S(n1157), .Y(n521) );
  MUX2X1 U2629 ( .B(n525), .A(n526), .S(n1157), .Y(n524) );
  MUX2X1 U2630 ( .B(n528), .A(n529), .S(n1157), .Y(n527) );
  MUX2X1 U2631 ( .B(n531), .A(n532), .S(n1191), .Y(n530) );
  MUX2X1 U2632 ( .B(n534), .A(n535), .S(n1157), .Y(n533) );
  MUX2X1 U2633 ( .B(n537), .A(n538), .S(n1157), .Y(n536) );
  MUX2X1 U2634 ( .B(n540), .A(n541), .S(n1157), .Y(n539) );
  MUX2X1 U2635 ( .B(n543), .A(n544), .S(n1157), .Y(n542) );
  MUX2X1 U2636 ( .B(n546), .A(n547), .S(n1191), .Y(n545) );
  MUX2X1 U2637 ( .B(n549), .A(n550), .S(n1157), .Y(n548) );
  MUX2X1 U2638 ( .B(n552), .A(n553), .S(n1157), .Y(n551) );
  MUX2X1 U2639 ( .B(n555), .A(n556), .S(n1157), .Y(n554) );
  MUX2X1 U2640 ( .B(n558), .A(n559), .S(n1157), .Y(n557) );
  MUX2X1 U2641 ( .B(n561), .A(n562), .S(n1191), .Y(n560) );
  MUX2X1 U2642 ( .B(n564), .A(n565), .S(n1158), .Y(n563) );
  MUX2X1 U2643 ( .B(n567), .A(n568), .S(n1158), .Y(n566) );
  MUX2X1 U2644 ( .B(n570), .A(n571), .S(n1158), .Y(n569) );
  MUX2X1 U2645 ( .B(n573), .A(n574), .S(n1158), .Y(n572) );
  MUX2X1 U2646 ( .B(n576), .A(n577), .S(n1191), .Y(n575) );
  MUX2X1 U2647 ( .B(n578), .A(n579), .S(n18), .Y(data_out[7]) );
  MUX2X1 U2648 ( .B(n581), .A(n582), .S(n1158), .Y(n580) );
  MUX2X1 U2649 ( .B(n584), .A(n585), .S(n1158), .Y(n583) );
  MUX2X1 U2650 ( .B(n587), .A(n588), .S(n1158), .Y(n586) );
  MUX2X1 U2651 ( .B(n590), .A(n591), .S(n1158), .Y(n589) );
  MUX2X1 U2652 ( .B(n593), .A(n594), .S(n1191), .Y(n592) );
  MUX2X1 U2653 ( .B(n596), .A(n597), .S(n1158), .Y(n595) );
  MUX2X1 U2654 ( .B(n599), .A(n600), .S(n1158), .Y(n598) );
  MUX2X1 U2655 ( .B(n602), .A(n603), .S(n1158), .Y(n601) );
  MUX2X1 U2656 ( .B(n605), .A(n606), .S(n1158), .Y(n604) );
  MUX2X1 U2657 ( .B(n608), .A(n609), .S(n1191), .Y(n607) );
  MUX2X1 U2658 ( .B(n611), .A(n612), .S(n1159), .Y(n610) );
  MUX2X1 U2659 ( .B(n614), .A(n615), .S(n1159), .Y(n613) );
  MUX2X1 U2660 ( .B(n617), .A(n618), .S(n1159), .Y(n616) );
  MUX2X1 U2661 ( .B(n620), .A(n621), .S(n1159), .Y(n619) );
  MUX2X1 U2662 ( .B(n623), .A(n624), .S(n1191), .Y(n622) );
  MUX2X1 U2663 ( .B(n626), .A(n627), .S(n1159), .Y(n625) );
  MUX2X1 U2664 ( .B(n629), .A(n630), .S(n1159), .Y(n628) );
  MUX2X1 U2665 ( .B(n632), .A(n633), .S(n1159), .Y(n631) );
  MUX2X1 U2666 ( .B(n635), .A(n636), .S(n1159), .Y(n634) );
  MUX2X1 U2667 ( .B(n638), .A(n639), .S(n1191), .Y(n637) );
  MUX2X1 U2668 ( .B(n640), .A(n641), .S(n18), .Y(data_out[8]) );
  MUX2X1 U2669 ( .B(n643), .A(n644), .S(n1159), .Y(n642) );
  MUX2X1 U2670 ( .B(n646), .A(n647), .S(n1159), .Y(n645) );
  MUX2X1 U2671 ( .B(n649), .A(n650), .S(n1159), .Y(n648) );
  MUX2X1 U2672 ( .B(n652), .A(n653), .S(n1159), .Y(n651) );
  MUX2X1 U2673 ( .B(n655), .A(n656), .S(n1191), .Y(n654) );
  MUX2X1 U2674 ( .B(n658), .A(n659), .S(n1160), .Y(n657) );
  MUX2X1 U2675 ( .B(n661), .A(n662), .S(n1160), .Y(n660) );
  MUX2X1 U2676 ( .B(n664), .A(n665), .S(n1160), .Y(n663) );
  MUX2X1 U2677 ( .B(n667), .A(n668), .S(n1160), .Y(n666) );
  MUX2X1 U2678 ( .B(n670), .A(n671), .S(n1191), .Y(n669) );
  MUX2X1 U2679 ( .B(n673), .A(n674), .S(n1160), .Y(n672) );
  MUX2X1 U2680 ( .B(n676), .A(n677), .S(n1160), .Y(n675) );
  MUX2X1 U2681 ( .B(n679), .A(n680), .S(n1160), .Y(n678) );
  MUX2X1 U2682 ( .B(n682), .A(n683), .S(n1160), .Y(n681) );
  MUX2X1 U2683 ( .B(n685), .A(n686), .S(n1191), .Y(n684) );
  MUX2X1 U2684 ( .B(n688), .A(n689), .S(n1160), .Y(n687) );
  MUX2X1 U2685 ( .B(n691), .A(n692), .S(n1160), .Y(n690) );
  MUX2X1 U2686 ( .B(n694), .A(n695), .S(n1160), .Y(n693) );
  MUX2X1 U2687 ( .B(n697), .A(n698), .S(n1160), .Y(n696) );
  MUX2X1 U2688 ( .B(n700), .A(n701), .S(n1191), .Y(n699) );
  MUX2X1 U2689 ( .B(n702), .A(n703), .S(n18), .Y(data_out[9]) );
  MUX2X1 U2690 ( .B(n705), .A(n706), .S(n1161), .Y(n704) );
  MUX2X1 U2691 ( .B(n708), .A(n709), .S(n1161), .Y(n707) );
  MUX2X1 U2692 ( .B(n711), .A(n712), .S(n1161), .Y(n710) );
  MUX2X1 U2693 ( .B(n714), .A(n715), .S(n1161), .Y(n713) );
  MUX2X1 U2694 ( .B(n717), .A(n718), .S(n1192), .Y(n716) );
  MUX2X1 U2695 ( .B(n720), .A(n721), .S(n1161), .Y(n719) );
  MUX2X1 U2696 ( .B(n723), .A(n724), .S(n1161), .Y(n722) );
  MUX2X1 U2697 ( .B(n726), .A(n727), .S(n1161), .Y(n725) );
  MUX2X1 U2698 ( .B(n729), .A(n730), .S(n1161), .Y(n728) );
  MUX2X1 U2699 ( .B(n732), .A(n733), .S(n1192), .Y(n731) );
  MUX2X1 U2700 ( .B(n735), .A(n736), .S(n1161), .Y(n734) );
  MUX2X1 U2701 ( .B(n738), .A(n739), .S(n1161), .Y(n737) );
  MUX2X1 U2702 ( .B(n741), .A(n742), .S(n1161), .Y(n740) );
  MUX2X1 U2703 ( .B(n744), .A(n745), .S(n1161), .Y(n743) );
  MUX2X1 U2704 ( .B(n747), .A(n748), .S(n1192), .Y(n746) );
  MUX2X1 U2705 ( .B(n750), .A(n751), .S(n1162), .Y(n749) );
  MUX2X1 U2706 ( .B(n753), .A(n754), .S(n1162), .Y(n752) );
  MUX2X1 U2707 ( .B(n756), .A(n757), .S(n1162), .Y(n755) );
  MUX2X1 U2708 ( .B(n759), .A(n760), .S(n1162), .Y(n758) );
  MUX2X1 U2709 ( .B(n762), .A(n763), .S(n1192), .Y(n761) );
  MUX2X1 U2710 ( .B(n764), .A(n765), .S(n18), .Y(data_out[10]) );
  MUX2X1 U2711 ( .B(n767), .A(n768), .S(n1162), .Y(n766) );
  MUX2X1 U2712 ( .B(n770), .A(n771), .S(n1162), .Y(n769) );
  MUX2X1 U2713 ( .B(n773), .A(n774), .S(n1162), .Y(n772) );
  MUX2X1 U2714 ( .B(n776), .A(n777), .S(n1162), .Y(n775) );
  MUX2X1 U2715 ( .B(n779), .A(n780), .S(n1192), .Y(n778) );
  MUX2X1 U2716 ( .B(n782), .A(n783), .S(n1162), .Y(n781) );
  MUX2X1 U2717 ( .B(n785), .A(n786), .S(n1162), .Y(n784) );
  MUX2X1 U2718 ( .B(n788), .A(n789), .S(n1162), .Y(n787) );
  MUX2X1 U2719 ( .B(n791), .A(n792), .S(n1162), .Y(n790) );
  MUX2X1 U2720 ( .B(n794), .A(n795), .S(n1192), .Y(n793) );
  MUX2X1 U2721 ( .B(n797), .A(n798), .S(n1163), .Y(n796) );
  MUX2X1 U2722 ( .B(n800), .A(n801), .S(n1163), .Y(n799) );
  MUX2X1 U2723 ( .B(n803), .A(n804), .S(n1163), .Y(n802) );
  MUX2X1 U2724 ( .B(n806), .A(n807), .S(n1163), .Y(n805) );
  MUX2X1 U2725 ( .B(n809), .A(n810), .S(n1192), .Y(n808) );
  MUX2X1 U2726 ( .B(n812), .A(n813), .S(n1163), .Y(n811) );
  MUX2X1 U2727 ( .B(n815), .A(n816), .S(n1163), .Y(n814) );
  MUX2X1 U2728 ( .B(n818), .A(n819), .S(n1163), .Y(n817) );
  MUX2X1 U2729 ( .B(n821), .A(n822), .S(n1163), .Y(n820) );
  MUX2X1 U2730 ( .B(n824), .A(n825), .S(n1192), .Y(n823) );
  MUX2X1 U2731 ( .B(n826), .A(n827), .S(n18), .Y(data_out[11]) );
  MUX2X1 U2732 ( .B(n829), .A(n830), .S(n1163), .Y(n828) );
  MUX2X1 U2733 ( .B(n832), .A(n833), .S(n1163), .Y(n831) );
  MUX2X1 U2734 ( .B(n835), .A(n836), .S(n1163), .Y(n834) );
  MUX2X1 U2735 ( .B(n838), .A(n839), .S(n1163), .Y(n837) );
  MUX2X1 U2736 ( .B(n841), .A(n842), .S(n1192), .Y(n840) );
  MUX2X1 U2737 ( .B(n844), .A(n845), .S(n1164), .Y(n843) );
  MUX2X1 U2738 ( .B(n847), .A(n848), .S(n1164), .Y(n846) );
  MUX2X1 U2739 ( .B(n850), .A(n851), .S(n1164), .Y(n849) );
  MUX2X1 U2740 ( .B(n853), .A(n854), .S(n1164), .Y(n852) );
  MUX2X1 U2741 ( .B(n856), .A(n857), .S(n1192), .Y(n855) );
  MUX2X1 U2742 ( .B(n859), .A(n860), .S(n1164), .Y(n858) );
  MUX2X1 U2743 ( .B(n862), .A(n863), .S(n1164), .Y(n861) );
  MUX2X1 U2744 ( .B(n865), .A(n866), .S(n1164), .Y(n864) );
  MUX2X1 U2745 ( .B(n868), .A(n869), .S(n1164), .Y(n867) );
  MUX2X1 U2746 ( .B(n871), .A(n872), .S(n1192), .Y(n870) );
  MUX2X1 U2747 ( .B(n874), .A(n875), .S(n1164), .Y(n873) );
  MUX2X1 U2748 ( .B(n877), .A(n878), .S(n1164), .Y(n876) );
  MUX2X1 U2749 ( .B(n880), .A(n881), .S(n1164), .Y(n879) );
  MUX2X1 U2750 ( .B(n883), .A(n884), .S(n1164), .Y(n882) );
  MUX2X1 U2751 ( .B(n886), .A(n887), .S(n1192), .Y(n885) );
  MUX2X1 U2752 ( .B(n888), .A(n889), .S(n18), .Y(data_out[12]) );
  MUX2X1 U2753 ( .B(n891), .A(n892), .S(n1165), .Y(n890) );
  MUX2X1 U2754 ( .B(n894), .A(n895), .S(n1165), .Y(n893) );
  MUX2X1 U2755 ( .B(n897), .A(n898), .S(n1165), .Y(n896) );
  MUX2X1 U2756 ( .B(n900), .A(n901), .S(n1165), .Y(n899) );
  MUX2X1 U2757 ( .B(n903), .A(n904), .S(n1193), .Y(n902) );
  MUX2X1 U2758 ( .B(n906), .A(n907), .S(n1165), .Y(n905) );
  MUX2X1 U2759 ( .B(n909), .A(n910), .S(n1165), .Y(n908) );
  MUX2X1 U2760 ( .B(n912), .A(n913), .S(n1165), .Y(n911) );
  MUX2X1 U2761 ( .B(n915), .A(n916), .S(n1165), .Y(n914) );
  MUX2X1 U2762 ( .B(n918), .A(n919), .S(n1193), .Y(n917) );
  MUX2X1 U2763 ( .B(n921), .A(n922), .S(n1165), .Y(n920) );
  MUX2X1 U2764 ( .B(n924), .A(n925), .S(n1165), .Y(n923) );
  MUX2X1 U2765 ( .B(n927), .A(n928), .S(n1165), .Y(n926) );
  MUX2X1 U2766 ( .B(n930), .A(n931), .S(n1165), .Y(n929) );
  MUX2X1 U2767 ( .B(n933), .A(n934), .S(n1193), .Y(n932) );
  MUX2X1 U2768 ( .B(n936), .A(n937), .S(n1166), .Y(n935) );
  MUX2X1 U2769 ( .B(n939), .A(n940), .S(n1166), .Y(n938) );
  MUX2X1 U2770 ( .B(n942), .A(n943), .S(n1166), .Y(n941) );
  MUX2X1 U2771 ( .B(n945), .A(n946), .S(n1166), .Y(n944) );
  MUX2X1 U2772 ( .B(n948), .A(n949), .S(n1193), .Y(n947) );
  MUX2X1 U2773 ( .B(n950), .A(n951), .S(n18), .Y(data_out[13]) );
  MUX2X1 U2774 ( .B(n953), .A(n954), .S(n1166), .Y(n952) );
  MUX2X1 U2775 ( .B(n956), .A(n957), .S(n1166), .Y(n955) );
  MUX2X1 U2776 ( .B(n959), .A(n960), .S(n1166), .Y(n958) );
  MUX2X1 U2777 ( .B(n962), .A(n963), .S(n1166), .Y(n961) );
  MUX2X1 U2778 ( .B(n965), .A(n966), .S(n1193), .Y(n964) );
  MUX2X1 U2779 ( .B(n968), .A(n969), .S(n1166), .Y(n967) );
  MUX2X1 U2780 ( .B(n971), .A(n972), .S(n1166), .Y(n970) );
  MUX2X1 U2781 ( .B(n974), .A(n975), .S(n1166), .Y(n973) );
  MUX2X1 U2782 ( .B(n977), .A(n978), .S(n1166), .Y(n976) );
  MUX2X1 U2783 ( .B(n980), .A(n981), .S(n1193), .Y(n979) );
  MUX2X1 U2784 ( .B(n983), .A(n984), .S(n1167), .Y(n982) );
  MUX2X1 U2785 ( .B(n986), .A(n987), .S(n1167), .Y(n985) );
  MUX2X1 U2786 ( .B(n989), .A(n990), .S(n1167), .Y(n988) );
  MUX2X1 U2787 ( .B(n992), .A(n993), .S(n1167), .Y(n991) );
  MUX2X1 U2788 ( .B(n995), .A(n996), .S(n1193), .Y(n994) );
  MUX2X1 U2789 ( .B(n998), .A(n999), .S(n1167), .Y(n997) );
  MUX2X1 U2790 ( .B(n1001), .A(n1002), .S(n1167), .Y(n1000) );
  MUX2X1 U2791 ( .B(n1004), .A(n1005), .S(n1167), .Y(n1003) );
  MUX2X1 U2792 ( .B(n1007), .A(n1008), .S(n1167), .Y(n1006) );
  MUX2X1 U2793 ( .B(n1010), .A(n1011), .S(n1193), .Y(n1009) );
  MUX2X1 U2794 ( .B(n1012), .A(n1013), .S(n18), .Y(data_out[14]) );
  MUX2X1 U2795 ( .B(n1015), .A(n1016), .S(n1167), .Y(n1014) );
  MUX2X1 U2796 ( .B(n1018), .A(n1019), .S(n1167), .Y(n1017) );
  MUX2X1 U2797 ( .B(n1021), .A(n1022), .S(n1167), .Y(n1020) );
  MUX2X1 U2798 ( .B(n1024), .A(n1025), .S(n1167), .Y(n1023) );
  MUX2X1 U2799 ( .B(n1027), .A(n1028), .S(n1193), .Y(n1026) );
  MUX2X1 U2800 ( .B(n1030), .A(n1031), .S(n1168), .Y(n1029) );
  MUX2X1 U2801 ( .B(n1033), .A(n1034), .S(n1168), .Y(n1032) );
  MUX2X1 U2802 ( .B(n1036), .A(n1037), .S(n1168), .Y(n1035) );
  MUX2X1 U2803 ( .B(n1039), .A(n1040), .S(n1168), .Y(n1038) );
  MUX2X1 U2804 ( .B(n1042), .A(n1043), .S(n1193), .Y(n1041) );
  MUX2X1 U2805 ( .B(n1045), .A(n1046), .S(n1168), .Y(n1044) );
  MUX2X1 U2806 ( .B(n1048), .A(n1049), .S(n1168), .Y(n1047) );
  MUX2X1 U2807 ( .B(n1051), .A(n1052), .S(n1168), .Y(n1050) );
  MUX2X1 U2808 ( .B(n1054), .A(n1055), .S(n1168), .Y(n1053) );
  MUX2X1 U2809 ( .B(n1057), .A(n1058), .S(n1193), .Y(n1056) );
  MUX2X1 U2810 ( .B(n1060), .A(n1061), .S(n1168), .Y(n1059) );
  MUX2X1 U2811 ( .B(n1063), .A(n1064), .S(n1168), .Y(n1062) );
  MUX2X1 U2812 ( .B(n1066), .A(n1067), .S(n1168), .Y(n1065) );
  MUX2X1 U2813 ( .B(n1069), .A(n1070), .S(n1168), .Y(n1068) );
  MUX2X1 U2814 ( .B(n1072), .A(n1073), .S(n1193), .Y(n1071) );
  MUX2X1 U2815 ( .B(n1074), .A(n1075), .S(n18), .Y(data_out[15]) );
  MUX2X1 U2816 ( .B(arr[992]), .A(arr[1008]), .S(n1076), .Y(n73) );
  MUX2X1 U2817 ( .B(arr[960]), .A(arr[976]), .S(n1076), .Y(n72) );
  MUX2X1 U2818 ( .B(arr[928]), .A(arr[944]), .S(n1076), .Y(n76) );
  MUX2X1 U2819 ( .B(arr[896]), .A(arr[912]), .S(n1076), .Y(n75) );
  MUX2X1 U2820 ( .B(n74), .A(n71), .S(n1177), .Y(n85) );
  MUX2X1 U2821 ( .B(arr[864]), .A(arr[880]), .S(n1076), .Y(n79) );
  MUX2X1 U2822 ( .B(arr[832]), .A(arr[848]), .S(n1076), .Y(n78) );
  MUX2X1 U2823 ( .B(arr[800]), .A(arr[816]), .S(n1076), .Y(n82) );
  MUX2X1 U2824 ( .B(arr[768]), .A(arr[784]), .S(n1076), .Y(n81) );
  MUX2X1 U2825 ( .B(n80), .A(n77), .S(n1177), .Y(n84) );
  MUX2X1 U2826 ( .B(arr[736]), .A(arr[752]), .S(n1077), .Y(n101) );
  MUX2X1 U2827 ( .B(arr[704]), .A(arr[720]), .S(n1077), .Y(n100) );
  MUX2X1 U2828 ( .B(arr[672]), .A(arr[688]), .S(n1077), .Y(n104) );
  MUX2X1 U2829 ( .B(arr[640]), .A(arr[656]), .S(n1077), .Y(n103) );
  MUX2X1 U2830 ( .B(n102), .A(n99), .S(n1177), .Y(n113) );
  MUX2X1 U2831 ( .B(arr[608]), .A(arr[624]), .S(n1077), .Y(n107) );
  MUX2X1 U2832 ( .B(arr[576]), .A(arr[592]), .S(n1077), .Y(n106) );
  MUX2X1 U2833 ( .B(arr[544]), .A(arr[560]), .S(n1077), .Y(n110) );
  MUX2X1 U2834 ( .B(arr[512]), .A(arr[528]), .S(n1077), .Y(n109) );
  MUX2X1 U2835 ( .B(n108), .A(n105), .S(n1177), .Y(n112) );
  MUX2X1 U2836 ( .B(n111), .A(n83), .S(n17), .Y(n145) );
  MUX2X1 U2837 ( .B(arr[480]), .A(arr[496]), .S(n1077), .Y(n116) );
  MUX2X1 U2838 ( .B(arr[448]), .A(arr[464]), .S(n1077), .Y(n115) );
  MUX2X1 U2839 ( .B(arr[416]), .A(arr[432]), .S(n1077), .Y(n119) );
  MUX2X1 U2840 ( .B(arr[384]), .A(arr[400]), .S(n1077), .Y(n118) );
  MUX2X1 U2841 ( .B(n117), .A(n114), .S(n1177), .Y(n128) );
  MUX2X1 U2842 ( .B(arr[352]), .A(arr[368]), .S(n1078), .Y(n122) );
  MUX2X1 U2843 ( .B(arr[320]), .A(arr[336]), .S(n1078), .Y(n121) );
  MUX2X1 U2844 ( .B(arr[288]), .A(arr[304]), .S(n1078), .Y(n125) );
  MUX2X1 U2845 ( .B(arr[256]), .A(arr[272]), .S(n1078), .Y(n124) );
  MUX2X1 U2846 ( .B(n123), .A(n120), .S(n1177), .Y(n127) );
  MUX2X1 U2847 ( .B(arr[224]), .A(arr[240]), .S(n1078), .Y(n131) );
  MUX2X1 U2848 ( .B(arr[192]), .A(arr[208]), .S(n1078), .Y(n130) );
  MUX2X1 U2849 ( .B(arr[160]), .A(arr[176]), .S(n1078), .Y(n134) );
  MUX2X1 U2850 ( .B(arr[128]), .A(arr[144]), .S(n1078), .Y(n133) );
  MUX2X1 U2851 ( .B(n132), .A(n129), .S(n1177), .Y(n143) );
  MUX2X1 U2852 ( .B(arr[96]), .A(arr[112]), .S(n1078), .Y(n137) );
  MUX2X1 U2853 ( .B(arr[64]), .A(arr[80]), .S(n1078), .Y(n136) );
  MUX2X1 U2854 ( .B(arr[32]), .A(arr[48]), .S(n1078), .Y(n140) );
  MUX2X1 U2855 ( .B(arr[0]), .A(arr[16]), .S(n1078), .Y(n139) );
  MUX2X1 U2856 ( .B(n138), .A(n135), .S(n1177), .Y(n142) );
  MUX2X1 U2857 ( .B(n141), .A(n126), .S(n17), .Y(n144) );
  MUX2X1 U2858 ( .B(arr[993]), .A(arr[1009]), .S(n1079), .Y(n148) );
  MUX2X1 U2859 ( .B(arr[961]), .A(arr[977]), .S(n1079), .Y(n147) );
  MUX2X1 U2860 ( .B(arr[929]), .A(arr[945]), .S(n1079), .Y(n151) );
  MUX2X1 U2861 ( .B(arr[897]), .A(arr[913]), .S(n1079), .Y(n150) );
  MUX2X1 U2862 ( .B(n149), .A(n146), .S(n1178), .Y(n160) );
  MUX2X1 U2863 ( .B(arr[865]), .A(arr[881]), .S(n1079), .Y(n154) );
  MUX2X1 U2864 ( .B(arr[833]), .A(arr[849]), .S(n1079), .Y(n153) );
  MUX2X1 U2865 ( .B(arr[801]), .A(arr[817]), .S(n1079), .Y(n157) );
  MUX2X1 U2866 ( .B(arr[769]), .A(arr[785]), .S(n1079), .Y(n156) );
  MUX2X1 U2867 ( .B(n155), .A(n152), .S(n1178), .Y(n159) );
  MUX2X1 U2868 ( .B(arr[737]), .A(arr[753]), .S(n1079), .Y(n163) );
  MUX2X1 U2869 ( .B(arr[705]), .A(arr[721]), .S(n1079), .Y(n162) );
  MUX2X1 U2870 ( .B(arr[673]), .A(arr[689]), .S(n1079), .Y(n166) );
  MUX2X1 U2871 ( .B(arr[641]), .A(arr[657]), .S(n1079), .Y(n165) );
  MUX2X1 U2872 ( .B(n164), .A(n161), .S(n1178), .Y(n175) );
  MUX2X1 U2873 ( .B(arr[609]), .A(arr[625]), .S(n1080), .Y(n169) );
  MUX2X1 U2874 ( .B(arr[577]), .A(arr[593]), .S(n1080), .Y(n168) );
  MUX2X1 U2875 ( .B(arr[545]), .A(arr[561]), .S(n1080), .Y(n172) );
  MUX2X1 U2876 ( .B(arr[513]), .A(arr[529]), .S(n1080), .Y(n171) );
  MUX2X1 U2877 ( .B(n170), .A(n167), .S(n1178), .Y(n174) );
  MUX2X1 U2878 ( .B(n173), .A(n158), .S(n17), .Y(n207) );
  MUX2X1 U2879 ( .B(arr[481]), .A(arr[497]), .S(n1080), .Y(n178) );
  MUX2X1 U2880 ( .B(arr[449]), .A(arr[465]), .S(n1080), .Y(n177) );
  MUX2X1 U2881 ( .B(arr[417]), .A(arr[433]), .S(n1080), .Y(n181) );
  MUX2X1 U2882 ( .B(arr[385]), .A(arr[401]), .S(n1080), .Y(n180) );
  MUX2X1 U2883 ( .B(n179), .A(n176), .S(n1178), .Y(n190) );
  MUX2X1 U2884 ( .B(arr[353]), .A(arr[369]), .S(n1080), .Y(n184) );
  MUX2X1 U2885 ( .B(arr[321]), .A(arr[337]), .S(n1080), .Y(n183) );
  MUX2X1 U2886 ( .B(arr[289]), .A(arr[305]), .S(n1080), .Y(n187) );
  MUX2X1 U2887 ( .B(arr[257]), .A(arr[273]), .S(n1080), .Y(n186) );
  MUX2X1 U2888 ( .B(n185), .A(n182), .S(n1178), .Y(n189) );
  MUX2X1 U2889 ( .B(arr[225]), .A(arr[241]), .S(n1081), .Y(n193) );
  MUX2X1 U2890 ( .B(arr[193]), .A(arr[209]), .S(n1081), .Y(n192) );
  MUX2X1 U2891 ( .B(arr[161]), .A(arr[177]), .S(n1081), .Y(n196) );
  MUX2X1 U2892 ( .B(arr[129]), .A(arr[145]), .S(n1081), .Y(n195) );
  MUX2X1 U2893 ( .B(n194), .A(n191), .S(n1178), .Y(n205) );
  MUX2X1 U2894 ( .B(arr[97]), .A(arr[113]), .S(n1081), .Y(n199) );
  MUX2X1 U2895 ( .B(arr[65]), .A(arr[81]), .S(n1081), .Y(n198) );
  MUX2X1 U2896 ( .B(arr[33]), .A(arr[49]), .S(n1081), .Y(n202) );
  MUX2X1 U2897 ( .B(arr[1]), .A(arr[17]), .S(n1081), .Y(n201) );
  MUX2X1 U2898 ( .B(n200), .A(n197), .S(n1178), .Y(n204) );
  MUX2X1 U2899 ( .B(n203), .A(n188), .S(n17), .Y(n206) );
  MUX2X1 U2900 ( .B(arr[994]), .A(arr[1010]), .S(n1081), .Y(n210) );
  MUX2X1 U2901 ( .B(arr[962]), .A(arr[978]), .S(n1081), .Y(n209) );
  MUX2X1 U2902 ( .B(arr[930]), .A(arr[946]), .S(n1081), .Y(n213) );
  MUX2X1 U2903 ( .B(arr[898]), .A(arr[914]), .S(n1081), .Y(n212) );
  MUX2X1 U2904 ( .B(n211), .A(n208), .S(n1178), .Y(n222) );
  MUX2X1 U2905 ( .B(arr[866]), .A(arr[882]), .S(n1082), .Y(n216) );
  MUX2X1 U2906 ( .B(arr[834]), .A(arr[850]), .S(n1082), .Y(n215) );
  MUX2X1 U2907 ( .B(arr[802]), .A(arr[818]), .S(n1082), .Y(n219) );
  MUX2X1 U2908 ( .B(arr[770]), .A(arr[786]), .S(n1082), .Y(n218) );
  MUX2X1 U2909 ( .B(n217), .A(n214), .S(n1178), .Y(n221) );
  MUX2X1 U2910 ( .B(arr[738]), .A(arr[754]), .S(n1082), .Y(n225) );
  MUX2X1 U2911 ( .B(arr[706]), .A(arr[722]), .S(n1082), .Y(n224) );
  MUX2X1 U2912 ( .B(arr[674]), .A(arr[690]), .S(n1082), .Y(n228) );
  MUX2X1 U2913 ( .B(arr[642]), .A(arr[658]), .S(n1082), .Y(n227) );
  MUX2X1 U2914 ( .B(n226), .A(n223), .S(n1178), .Y(n237) );
  MUX2X1 U2915 ( .B(arr[610]), .A(arr[626]), .S(n1082), .Y(n231) );
  MUX2X1 U2916 ( .B(arr[578]), .A(arr[594]), .S(n1082), .Y(n230) );
  MUX2X1 U2917 ( .B(arr[546]), .A(arr[562]), .S(n1082), .Y(n234) );
  MUX2X1 U2918 ( .B(arr[514]), .A(arr[530]), .S(n1082), .Y(n233) );
  MUX2X1 U2919 ( .B(n232), .A(n229), .S(n1178), .Y(n236) );
  MUX2X1 U2920 ( .B(n235), .A(n220), .S(n17), .Y(n269) );
  MUX2X1 U2921 ( .B(arr[482]), .A(arr[498]), .S(n1083), .Y(n240) );
  MUX2X1 U2922 ( .B(arr[450]), .A(arr[466]), .S(n1083), .Y(n239) );
  MUX2X1 U2923 ( .B(arr[418]), .A(arr[434]), .S(n1083), .Y(n243) );
  MUX2X1 U2924 ( .B(arr[386]), .A(arr[402]), .S(n1083), .Y(n242) );
  MUX2X1 U2925 ( .B(n241), .A(n238), .S(n1179), .Y(n252) );
  MUX2X1 U2926 ( .B(arr[354]), .A(arr[370]), .S(n1083), .Y(n246) );
  MUX2X1 U2927 ( .B(arr[322]), .A(arr[338]), .S(n1083), .Y(n245) );
  MUX2X1 U2928 ( .B(arr[290]), .A(arr[306]), .S(n1083), .Y(n249) );
  MUX2X1 U2929 ( .B(arr[258]), .A(arr[274]), .S(n1083), .Y(n248) );
  MUX2X1 U2930 ( .B(n247), .A(n244), .S(n1179), .Y(n251) );
  MUX2X1 U2931 ( .B(arr[226]), .A(arr[242]), .S(n1083), .Y(n255) );
  MUX2X1 U2932 ( .B(arr[194]), .A(arr[210]), .S(n1083), .Y(n254) );
  MUX2X1 U2933 ( .B(arr[162]), .A(arr[178]), .S(n1083), .Y(n258) );
  MUX2X1 U2934 ( .B(arr[130]), .A(arr[146]), .S(n1083), .Y(n257) );
  MUX2X1 U2935 ( .B(n256), .A(n253), .S(n1179), .Y(n267) );
  MUX2X1 U2936 ( .B(arr[98]), .A(arr[114]), .S(n1084), .Y(n261) );
  MUX2X1 U2937 ( .B(arr[66]), .A(arr[82]), .S(n1084), .Y(n260) );
  MUX2X1 U2938 ( .B(arr[34]), .A(arr[50]), .S(n1084), .Y(n264) );
  MUX2X1 U2939 ( .B(arr[2]), .A(arr[18]), .S(n1084), .Y(n263) );
  MUX2X1 U2940 ( .B(n262), .A(n259), .S(n1179), .Y(n266) );
  MUX2X1 U2941 ( .B(n265), .A(n250), .S(n17), .Y(n268) );
  MUX2X1 U2942 ( .B(arr[995]), .A(arr[1011]), .S(n1084), .Y(n272) );
  MUX2X1 U2943 ( .B(arr[963]), .A(arr[979]), .S(n1084), .Y(n271) );
  MUX2X1 U2944 ( .B(arr[931]), .A(arr[947]), .S(n1084), .Y(n275) );
  MUX2X1 U2945 ( .B(arr[899]), .A(arr[915]), .S(n1084), .Y(n274) );
  MUX2X1 U2946 ( .B(n273), .A(n270), .S(n1179), .Y(n284) );
  MUX2X1 U2947 ( .B(arr[867]), .A(arr[883]), .S(n1084), .Y(n278) );
  MUX2X1 U2948 ( .B(arr[835]), .A(arr[851]), .S(n1084), .Y(n277) );
  MUX2X1 U2949 ( .B(arr[803]), .A(arr[819]), .S(n1084), .Y(n281) );
  MUX2X1 U2950 ( .B(arr[771]), .A(arr[787]), .S(n1084), .Y(n280) );
  MUX2X1 U2951 ( .B(n279), .A(n276), .S(n1179), .Y(n283) );
  MUX2X1 U2952 ( .B(arr[739]), .A(arr[755]), .S(n1085), .Y(n287) );
  MUX2X1 U2953 ( .B(arr[707]), .A(arr[723]), .S(n1085), .Y(n286) );
  MUX2X1 U2954 ( .B(arr[675]), .A(arr[691]), .S(n1085), .Y(n290) );
  MUX2X1 U2955 ( .B(arr[643]), .A(arr[659]), .S(n1085), .Y(n289) );
  MUX2X1 U2956 ( .B(n288), .A(n285), .S(n1179), .Y(n299) );
  MUX2X1 U2957 ( .B(arr[611]), .A(arr[627]), .S(n1085), .Y(n293) );
  MUX2X1 U2958 ( .B(arr[579]), .A(arr[595]), .S(n1085), .Y(n292) );
  MUX2X1 U2959 ( .B(arr[547]), .A(arr[563]), .S(n1085), .Y(n296) );
  MUX2X1 U2960 ( .B(arr[515]), .A(arr[531]), .S(n1085), .Y(n295) );
  MUX2X1 U2961 ( .B(n294), .A(n291), .S(n1179), .Y(n298) );
  MUX2X1 U2962 ( .B(n297), .A(n282), .S(n17), .Y(n331) );
  MUX2X1 U2963 ( .B(arr[483]), .A(arr[499]), .S(n1085), .Y(n302) );
  MUX2X1 U2964 ( .B(arr[451]), .A(arr[467]), .S(n1085), .Y(n301) );
  MUX2X1 U2965 ( .B(arr[419]), .A(arr[435]), .S(n1085), .Y(n305) );
  MUX2X1 U2966 ( .B(arr[387]), .A(arr[403]), .S(n1085), .Y(n304) );
  MUX2X1 U2967 ( .B(n303), .A(n300), .S(n1179), .Y(n314) );
  MUX2X1 U2968 ( .B(arr[355]), .A(arr[371]), .S(n1086), .Y(n308) );
  MUX2X1 U2969 ( .B(arr[323]), .A(arr[339]), .S(n1086), .Y(n307) );
  MUX2X1 U2970 ( .B(arr[291]), .A(arr[307]), .S(n1086), .Y(n311) );
  MUX2X1 U2971 ( .B(arr[259]), .A(arr[275]), .S(n1086), .Y(n310) );
  MUX2X1 U2972 ( .B(n309), .A(n306), .S(n1179), .Y(n313) );
  MUX2X1 U2973 ( .B(arr[227]), .A(arr[243]), .S(n1086), .Y(n317) );
  MUX2X1 U2974 ( .B(arr[195]), .A(arr[211]), .S(n1086), .Y(n316) );
  MUX2X1 U2975 ( .B(arr[163]), .A(arr[179]), .S(n1086), .Y(n320) );
  MUX2X1 U2976 ( .B(arr[131]), .A(arr[147]), .S(n1086), .Y(n319) );
  MUX2X1 U2977 ( .B(n318), .A(n315), .S(n1179), .Y(n329) );
  MUX2X1 U2978 ( .B(arr[99]), .A(arr[115]), .S(n1086), .Y(n323) );
  MUX2X1 U2979 ( .B(arr[67]), .A(arr[83]), .S(n1086), .Y(n322) );
  MUX2X1 U2980 ( .B(arr[35]), .A(arr[51]), .S(n1086), .Y(n326) );
  MUX2X1 U2981 ( .B(arr[3]), .A(arr[19]), .S(n1086), .Y(n325) );
  MUX2X1 U2982 ( .B(n324), .A(n321), .S(n1179), .Y(n328) );
  MUX2X1 U2983 ( .B(n327), .A(n312), .S(n17), .Y(n330) );
  MUX2X1 U2984 ( .B(arr[996]), .A(arr[1012]), .S(n1087), .Y(n334) );
  MUX2X1 U2985 ( .B(arr[964]), .A(arr[980]), .S(n1087), .Y(n333) );
  MUX2X1 U2986 ( .B(arr[932]), .A(arr[948]), .S(n1087), .Y(n337) );
  MUX2X1 U2987 ( .B(arr[900]), .A(arr[916]), .S(n1087), .Y(n336) );
  MUX2X1 U2988 ( .B(n335), .A(n332), .S(n1180), .Y(n346) );
  MUX2X1 U2989 ( .B(arr[868]), .A(arr[884]), .S(n1087), .Y(n340) );
  MUX2X1 U2990 ( .B(arr[836]), .A(arr[852]), .S(n1087), .Y(n339) );
  MUX2X1 U2991 ( .B(arr[804]), .A(arr[820]), .S(n1087), .Y(n343) );
  MUX2X1 U2992 ( .B(arr[772]), .A(arr[788]), .S(n1087), .Y(n342) );
  MUX2X1 U2993 ( .B(n341), .A(n338), .S(n1180), .Y(n345) );
  MUX2X1 U2994 ( .B(arr[740]), .A(arr[756]), .S(n1087), .Y(n349) );
  MUX2X1 U2995 ( .B(arr[708]), .A(arr[724]), .S(n1087), .Y(n348) );
  MUX2X1 U2996 ( .B(arr[676]), .A(arr[692]), .S(n1087), .Y(n352) );
  MUX2X1 U2997 ( .B(arr[644]), .A(arr[660]), .S(n1087), .Y(n351) );
  MUX2X1 U2998 ( .B(n350), .A(n347), .S(n1180), .Y(n361) );
  MUX2X1 U2999 ( .B(arr[612]), .A(arr[628]), .S(n1088), .Y(n355) );
  MUX2X1 U3000 ( .B(arr[580]), .A(arr[596]), .S(n1088), .Y(n354) );
  MUX2X1 U3001 ( .B(arr[548]), .A(arr[564]), .S(n1088), .Y(n358) );
  MUX2X1 U3002 ( .B(arr[516]), .A(arr[532]), .S(n1088), .Y(n357) );
  MUX2X1 U3003 ( .B(n356), .A(n353), .S(n1180), .Y(n360) );
  MUX2X1 U3004 ( .B(n359), .A(n344), .S(n17), .Y(n393) );
  MUX2X1 U3005 ( .B(arr[484]), .A(arr[500]), .S(n1088), .Y(n364) );
  MUX2X1 U3006 ( .B(arr[452]), .A(arr[468]), .S(n1088), .Y(n363) );
  MUX2X1 U3007 ( .B(arr[420]), .A(arr[436]), .S(n1088), .Y(n367) );
  MUX2X1 U3008 ( .B(arr[388]), .A(arr[404]), .S(n1088), .Y(n366) );
  MUX2X1 U3009 ( .B(n365), .A(n362), .S(n1180), .Y(n376) );
  MUX2X1 U3010 ( .B(arr[356]), .A(arr[372]), .S(n1088), .Y(n370) );
  MUX2X1 U3011 ( .B(arr[324]), .A(arr[340]), .S(n1088), .Y(n369) );
  MUX2X1 U3012 ( .B(arr[292]), .A(arr[308]), .S(n1088), .Y(n373) );
  MUX2X1 U3013 ( .B(arr[260]), .A(arr[276]), .S(n1088), .Y(n372) );
  MUX2X1 U3014 ( .B(n371), .A(n368), .S(n1180), .Y(n375) );
  MUX2X1 U3015 ( .B(arr[228]), .A(arr[244]), .S(n1089), .Y(n379) );
  MUX2X1 U3016 ( .B(arr[196]), .A(arr[212]), .S(n1089), .Y(n378) );
  MUX2X1 U3017 ( .B(arr[164]), .A(arr[180]), .S(n1089), .Y(n382) );
  MUX2X1 U3018 ( .B(arr[132]), .A(arr[148]), .S(n1089), .Y(n381) );
  MUX2X1 U3019 ( .B(n380), .A(n377), .S(n1180), .Y(n391) );
  MUX2X1 U3020 ( .B(arr[100]), .A(arr[116]), .S(n1089), .Y(n385) );
  MUX2X1 U3021 ( .B(arr[68]), .A(arr[84]), .S(n1089), .Y(n384) );
  MUX2X1 U3022 ( .B(arr[36]), .A(arr[52]), .S(n1089), .Y(n388) );
  MUX2X1 U3023 ( .B(arr[4]), .A(arr[20]), .S(n1089), .Y(n387) );
  MUX2X1 U3024 ( .B(n386), .A(n383), .S(n1180), .Y(n390) );
  MUX2X1 U3025 ( .B(n389), .A(n374), .S(n17), .Y(n392) );
  MUX2X1 U3026 ( .B(arr[997]), .A(arr[1013]), .S(n1089), .Y(n396) );
  MUX2X1 U3027 ( .B(arr[965]), .A(arr[981]), .S(n1089), .Y(n395) );
  MUX2X1 U3028 ( .B(arr[933]), .A(arr[949]), .S(n1089), .Y(n399) );
  MUX2X1 U3029 ( .B(arr[901]), .A(arr[917]), .S(n1089), .Y(n398) );
  MUX2X1 U3030 ( .B(n397), .A(n394), .S(n1180), .Y(n408) );
  MUX2X1 U3031 ( .B(arr[869]), .A(arr[885]), .S(n1090), .Y(n402) );
  MUX2X1 U3032 ( .B(arr[837]), .A(arr[853]), .S(n1090), .Y(n401) );
  MUX2X1 U3033 ( .B(arr[805]), .A(arr[821]), .S(n1090), .Y(n405) );
  MUX2X1 U3034 ( .B(arr[773]), .A(arr[789]), .S(n1090), .Y(n404) );
  MUX2X1 U3035 ( .B(n403), .A(n400), .S(n1180), .Y(n407) );
  MUX2X1 U3036 ( .B(arr[741]), .A(arr[757]), .S(n1090), .Y(n411) );
  MUX2X1 U3037 ( .B(arr[709]), .A(arr[725]), .S(n1090), .Y(n410) );
  MUX2X1 U3038 ( .B(arr[677]), .A(arr[693]), .S(n1090), .Y(n414) );
  MUX2X1 U3039 ( .B(arr[645]), .A(arr[661]), .S(n1090), .Y(n413) );
  MUX2X1 U3040 ( .B(n412), .A(n409), .S(n1180), .Y(n423) );
  MUX2X1 U3041 ( .B(arr[613]), .A(arr[629]), .S(n1090), .Y(n417) );
  MUX2X1 U3042 ( .B(arr[581]), .A(arr[597]), .S(n1090), .Y(n416) );
  MUX2X1 U3043 ( .B(arr[549]), .A(arr[565]), .S(n1090), .Y(n420) );
  MUX2X1 U3044 ( .B(arr[517]), .A(arr[533]), .S(n1090), .Y(n419) );
  MUX2X1 U3045 ( .B(n418), .A(n415), .S(n1180), .Y(n422) );
  MUX2X1 U3046 ( .B(n421), .A(n406), .S(n17), .Y(n455) );
  MUX2X1 U3047 ( .B(arr[485]), .A(arr[501]), .S(n1091), .Y(n426) );
  MUX2X1 U3048 ( .B(arr[453]), .A(arr[469]), .S(n1091), .Y(n425) );
  MUX2X1 U3049 ( .B(arr[421]), .A(arr[437]), .S(n1091), .Y(n429) );
  MUX2X1 U3050 ( .B(arr[389]), .A(arr[405]), .S(n1091), .Y(n428) );
  MUX2X1 U3051 ( .B(n427), .A(n424), .S(n1181), .Y(n438) );
  MUX2X1 U3052 ( .B(arr[357]), .A(arr[373]), .S(n1091), .Y(n432) );
  MUX2X1 U3053 ( .B(arr[325]), .A(arr[341]), .S(n1091), .Y(n431) );
  MUX2X1 U3054 ( .B(arr[293]), .A(arr[309]), .S(n1091), .Y(n435) );
  MUX2X1 U3055 ( .B(arr[261]), .A(arr[277]), .S(n1091), .Y(n434) );
  MUX2X1 U3056 ( .B(n433), .A(n430), .S(n1181), .Y(n437) );
  MUX2X1 U3057 ( .B(arr[229]), .A(arr[245]), .S(n1091), .Y(n441) );
  MUX2X1 U3058 ( .B(arr[197]), .A(arr[213]), .S(n1091), .Y(n440) );
  MUX2X1 U3059 ( .B(arr[165]), .A(arr[181]), .S(n1091), .Y(n444) );
  MUX2X1 U3060 ( .B(arr[133]), .A(arr[149]), .S(n1091), .Y(n443) );
  MUX2X1 U3061 ( .B(n442), .A(n439), .S(n1181), .Y(n453) );
  MUX2X1 U3062 ( .B(arr[101]), .A(arr[117]), .S(n1092), .Y(n447) );
  MUX2X1 U3063 ( .B(arr[69]), .A(arr[85]), .S(n1092), .Y(n446) );
  MUX2X1 U3064 ( .B(arr[37]), .A(arr[53]), .S(n1092), .Y(n450) );
  MUX2X1 U3065 ( .B(arr[5]), .A(arr[21]), .S(n1092), .Y(n449) );
  MUX2X1 U3066 ( .B(n448), .A(n445), .S(n1181), .Y(n452) );
  MUX2X1 U3067 ( .B(n451), .A(n436), .S(n17), .Y(n454) );
  MUX2X1 U3068 ( .B(arr[998]), .A(arr[1014]), .S(n1092), .Y(n458) );
  MUX2X1 U3069 ( .B(arr[966]), .A(arr[982]), .S(n1092), .Y(n457) );
  MUX2X1 U3070 ( .B(arr[934]), .A(arr[950]), .S(n1092), .Y(n461) );
  MUX2X1 U3071 ( .B(arr[902]), .A(arr[918]), .S(n1092), .Y(n460) );
  MUX2X1 U3072 ( .B(n459), .A(n456), .S(n1181), .Y(n470) );
  MUX2X1 U3073 ( .B(arr[870]), .A(arr[886]), .S(n1092), .Y(n464) );
  MUX2X1 U3074 ( .B(arr[838]), .A(arr[854]), .S(n1092), .Y(n463) );
  MUX2X1 U3075 ( .B(arr[806]), .A(arr[822]), .S(n1092), .Y(n467) );
  MUX2X1 U3076 ( .B(arr[774]), .A(arr[790]), .S(n1092), .Y(n466) );
  MUX2X1 U3077 ( .B(n465), .A(n462), .S(n1181), .Y(n469) );
  MUX2X1 U3078 ( .B(arr[742]), .A(arr[758]), .S(n1093), .Y(n473) );
  MUX2X1 U3079 ( .B(arr[710]), .A(arr[726]), .S(n1093), .Y(n472) );
  MUX2X1 U3080 ( .B(arr[678]), .A(arr[694]), .S(n1093), .Y(n476) );
  MUX2X1 U3081 ( .B(arr[646]), .A(arr[662]), .S(n1093), .Y(n475) );
  MUX2X1 U3082 ( .B(n474), .A(n471), .S(n1181), .Y(n485) );
  MUX2X1 U3083 ( .B(arr[614]), .A(arr[630]), .S(n1093), .Y(n479) );
  MUX2X1 U3084 ( .B(arr[582]), .A(arr[598]), .S(n1093), .Y(n478) );
  MUX2X1 U3085 ( .B(arr[550]), .A(arr[566]), .S(n1093), .Y(n482) );
  MUX2X1 U3086 ( .B(arr[518]), .A(arr[534]), .S(n1093), .Y(n481) );
  MUX2X1 U3087 ( .B(n480), .A(n477), .S(n1181), .Y(n484) );
  MUX2X1 U3088 ( .B(n483), .A(n468), .S(n17), .Y(n517) );
  MUX2X1 U3089 ( .B(arr[486]), .A(arr[502]), .S(n1093), .Y(n488) );
  MUX2X1 U3090 ( .B(arr[454]), .A(arr[470]), .S(n1093), .Y(n487) );
  MUX2X1 U3091 ( .B(arr[422]), .A(arr[438]), .S(n1093), .Y(n491) );
  MUX2X1 U3092 ( .B(arr[390]), .A(arr[406]), .S(n1093), .Y(n490) );
  MUX2X1 U3093 ( .B(n489), .A(n486), .S(n1181), .Y(n500) );
  MUX2X1 U3094 ( .B(arr[358]), .A(arr[374]), .S(n1094), .Y(n494) );
  MUX2X1 U3095 ( .B(arr[326]), .A(arr[342]), .S(n1094), .Y(n493) );
  MUX2X1 U3096 ( .B(arr[294]), .A(arr[310]), .S(n1094), .Y(n497) );
  MUX2X1 U3097 ( .B(arr[262]), .A(arr[278]), .S(n1094), .Y(n496) );
  MUX2X1 U3098 ( .B(n495), .A(n492), .S(n1181), .Y(n499) );
  MUX2X1 U3099 ( .B(arr[230]), .A(arr[246]), .S(n1094), .Y(n503) );
  MUX2X1 U3100 ( .B(arr[198]), .A(arr[214]), .S(n1094), .Y(n502) );
  MUX2X1 U3101 ( .B(arr[166]), .A(arr[182]), .S(n1094), .Y(n506) );
  MUX2X1 U3102 ( .B(arr[134]), .A(arr[150]), .S(n1094), .Y(n505) );
  MUX2X1 U3103 ( .B(n504), .A(n501), .S(n1181), .Y(n515) );
  MUX2X1 U3104 ( .B(arr[102]), .A(arr[118]), .S(n1094), .Y(n509) );
  MUX2X1 U3105 ( .B(arr[70]), .A(arr[86]), .S(n1094), .Y(n508) );
  MUX2X1 U3106 ( .B(arr[38]), .A(arr[54]), .S(n1094), .Y(n512) );
  MUX2X1 U3107 ( .B(arr[6]), .A(arr[22]), .S(n1094), .Y(n511) );
  MUX2X1 U3108 ( .B(n510), .A(n507), .S(n1181), .Y(n514) );
  MUX2X1 U3109 ( .B(n513), .A(n498), .S(n17), .Y(n516) );
  MUX2X1 U3110 ( .B(arr[999]), .A(arr[1015]), .S(n1095), .Y(n520) );
  MUX2X1 U3111 ( .B(arr[967]), .A(arr[983]), .S(n1095), .Y(n519) );
  MUX2X1 U3112 ( .B(arr[935]), .A(arr[951]), .S(n1095), .Y(n523) );
  MUX2X1 U3113 ( .B(arr[903]), .A(arr[919]), .S(n1095), .Y(n522) );
  MUX2X1 U3114 ( .B(n521), .A(n518), .S(n1182), .Y(n532) );
  MUX2X1 U3115 ( .B(arr[871]), .A(arr[887]), .S(n1095), .Y(n526) );
  MUX2X1 U3116 ( .B(arr[839]), .A(arr[855]), .S(n1095), .Y(n525) );
  MUX2X1 U3117 ( .B(arr[807]), .A(arr[823]), .S(n1095), .Y(n529) );
  MUX2X1 U3118 ( .B(arr[775]), .A(arr[791]), .S(n1095), .Y(n528) );
  MUX2X1 U3119 ( .B(n527), .A(n524), .S(n1182), .Y(n531) );
  MUX2X1 U3120 ( .B(arr[743]), .A(arr[759]), .S(n1095), .Y(n535) );
  MUX2X1 U3121 ( .B(arr[711]), .A(arr[727]), .S(n1095), .Y(n534) );
  MUX2X1 U3122 ( .B(arr[679]), .A(arr[695]), .S(n1095), .Y(n538) );
  MUX2X1 U3123 ( .B(arr[647]), .A(arr[663]), .S(n1095), .Y(n537) );
  MUX2X1 U3124 ( .B(n536), .A(n533), .S(n1182), .Y(n547) );
  MUX2X1 U3125 ( .B(arr[615]), .A(arr[631]), .S(n1096), .Y(n541) );
  MUX2X1 U3126 ( .B(arr[583]), .A(arr[599]), .S(n1096), .Y(n540) );
  MUX2X1 U3127 ( .B(arr[551]), .A(arr[567]), .S(n1096), .Y(n544) );
  MUX2X1 U3128 ( .B(arr[519]), .A(arr[535]), .S(n1096), .Y(n543) );
  MUX2X1 U3129 ( .B(n542), .A(n539), .S(n1182), .Y(n546) );
  MUX2X1 U3130 ( .B(n545), .A(n530), .S(n17), .Y(n579) );
  MUX2X1 U3131 ( .B(arr[487]), .A(arr[503]), .S(n1096), .Y(n550) );
  MUX2X1 U3132 ( .B(arr[455]), .A(arr[471]), .S(n1096), .Y(n549) );
  MUX2X1 U3133 ( .B(arr[423]), .A(arr[439]), .S(n1096), .Y(n553) );
  MUX2X1 U3134 ( .B(arr[391]), .A(arr[407]), .S(n1096), .Y(n552) );
  MUX2X1 U3135 ( .B(n551), .A(n548), .S(n1182), .Y(n562) );
  MUX2X1 U3136 ( .B(arr[359]), .A(arr[375]), .S(n1096), .Y(n556) );
  MUX2X1 U3137 ( .B(arr[327]), .A(arr[343]), .S(n1096), .Y(n555) );
  MUX2X1 U3138 ( .B(arr[295]), .A(arr[311]), .S(n1096), .Y(n559) );
  MUX2X1 U3139 ( .B(arr[263]), .A(arr[279]), .S(n1096), .Y(n558) );
  MUX2X1 U3140 ( .B(n557), .A(n554), .S(n1182), .Y(n561) );
  MUX2X1 U3141 ( .B(arr[231]), .A(arr[247]), .S(n1097), .Y(n565) );
  MUX2X1 U3142 ( .B(arr[199]), .A(arr[215]), .S(n1097), .Y(n564) );
  MUX2X1 U3143 ( .B(arr[167]), .A(arr[183]), .S(n1097), .Y(n568) );
  MUX2X1 U3144 ( .B(arr[135]), .A(arr[151]), .S(n1097), .Y(n567) );
  MUX2X1 U3145 ( .B(n566), .A(n563), .S(n1182), .Y(n577) );
  MUX2X1 U3146 ( .B(arr[103]), .A(arr[119]), .S(n1097), .Y(n571) );
  MUX2X1 U3147 ( .B(arr[71]), .A(arr[87]), .S(n1097), .Y(n570) );
  MUX2X1 U3148 ( .B(arr[39]), .A(arr[55]), .S(n1097), .Y(n574) );
  MUX2X1 U3149 ( .B(arr[7]), .A(arr[23]), .S(n1097), .Y(n573) );
  MUX2X1 U3150 ( .B(n572), .A(n569), .S(n1182), .Y(n576) );
  MUX2X1 U3151 ( .B(n575), .A(n560), .S(n17), .Y(n578) );
  MUX2X1 U3152 ( .B(arr[1000]), .A(arr[1016]), .S(n1097), .Y(n582) );
  MUX2X1 U3153 ( .B(arr[968]), .A(arr[984]), .S(n1097), .Y(n581) );
  MUX2X1 U3154 ( .B(arr[936]), .A(arr[952]), .S(n1097), .Y(n585) );
  MUX2X1 U3155 ( .B(arr[904]), .A(arr[920]), .S(n1097), .Y(n584) );
  MUX2X1 U3156 ( .B(n583), .A(n580), .S(n1182), .Y(n594) );
  MUX2X1 U3157 ( .B(arr[872]), .A(arr[888]), .S(n1098), .Y(n588) );
  MUX2X1 U3158 ( .B(arr[840]), .A(arr[856]), .S(n1098), .Y(n587) );
  MUX2X1 U3159 ( .B(arr[808]), .A(arr[824]), .S(n1098), .Y(n591) );
  MUX2X1 U3160 ( .B(arr[776]), .A(arr[792]), .S(n1098), .Y(n590) );
  MUX2X1 U3161 ( .B(n589), .A(n586), .S(n1182), .Y(n593) );
  MUX2X1 U3162 ( .B(arr[744]), .A(arr[760]), .S(n1098), .Y(n597) );
  MUX2X1 U3163 ( .B(arr[712]), .A(arr[728]), .S(n1098), .Y(n596) );
  MUX2X1 U3164 ( .B(arr[680]), .A(arr[696]), .S(n1098), .Y(n600) );
  MUX2X1 U3165 ( .B(arr[648]), .A(arr[664]), .S(n1098), .Y(n599) );
  MUX2X1 U3166 ( .B(n598), .A(n595), .S(n1182), .Y(n609) );
  MUX2X1 U3167 ( .B(arr[616]), .A(arr[632]), .S(n1098), .Y(n603) );
  MUX2X1 U3168 ( .B(arr[584]), .A(arr[600]), .S(n1098), .Y(n602) );
  MUX2X1 U3169 ( .B(arr[552]), .A(arr[568]), .S(n1098), .Y(n606) );
  MUX2X1 U3170 ( .B(arr[520]), .A(arr[536]), .S(n1098), .Y(n605) );
  MUX2X1 U3171 ( .B(n604), .A(n601), .S(n1182), .Y(n608) );
  MUX2X1 U3172 ( .B(n607), .A(n592), .S(n17), .Y(n641) );
  MUX2X1 U3173 ( .B(arr[488]), .A(arr[504]), .S(n1099), .Y(n612) );
  MUX2X1 U3174 ( .B(arr[456]), .A(arr[472]), .S(n1099), .Y(n611) );
  MUX2X1 U3175 ( .B(arr[424]), .A(arr[440]), .S(n1099), .Y(n615) );
  MUX2X1 U3176 ( .B(arr[392]), .A(arr[408]), .S(n1099), .Y(n614) );
  MUX2X1 U3177 ( .B(n613), .A(n610), .S(n1183), .Y(n624) );
  MUX2X1 U3178 ( .B(arr[360]), .A(arr[376]), .S(n1099), .Y(n618) );
  MUX2X1 U3179 ( .B(arr[328]), .A(arr[344]), .S(n1099), .Y(n617) );
  MUX2X1 U3180 ( .B(arr[296]), .A(arr[312]), .S(n1099), .Y(n621) );
  MUX2X1 U3181 ( .B(arr[264]), .A(arr[280]), .S(n1099), .Y(n620) );
  MUX2X1 U3182 ( .B(n619), .A(n616), .S(n1183), .Y(n623) );
  MUX2X1 U3183 ( .B(arr[232]), .A(arr[248]), .S(n1099), .Y(n627) );
  MUX2X1 U3184 ( .B(arr[200]), .A(arr[216]), .S(n1099), .Y(n626) );
  MUX2X1 U3185 ( .B(arr[168]), .A(arr[184]), .S(n1099), .Y(n630) );
  MUX2X1 U3186 ( .B(arr[136]), .A(arr[152]), .S(n1099), .Y(n629) );
  MUX2X1 U3187 ( .B(n628), .A(n625), .S(n1183), .Y(n639) );
  MUX2X1 U3188 ( .B(arr[104]), .A(arr[120]), .S(n1100), .Y(n633) );
  MUX2X1 U3189 ( .B(arr[72]), .A(arr[88]), .S(n1100), .Y(n632) );
  MUX2X1 U3190 ( .B(arr[40]), .A(arr[56]), .S(n1100), .Y(n636) );
  MUX2X1 U3191 ( .B(arr[8]), .A(arr[24]), .S(n1100), .Y(n635) );
  MUX2X1 U3192 ( .B(n634), .A(n631), .S(n1183), .Y(n638) );
  MUX2X1 U3193 ( .B(n637), .A(n622), .S(n17), .Y(n640) );
  MUX2X1 U3194 ( .B(arr[1001]), .A(arr[1017]), .S(n1100), .Y(n644) );
  MUX2X1 U3195 ( .B(arr[969]), .A(arr[985]), .S(n1100), .Y(n643) );
  MUX2X1 U3196 ( .B(arr[937]), .A(arr[953]), .S(n1100), .Y(n647) );
  MUX2X1 U3197 ( .B(arr[905]), .A(arr[921]), .S(n1100), .Y(n646) );
  MUX2X1 U3198 ( .B(n645), .A(n642), .S(n1183), .Y(n656) );
  MUX2X1 U3199 ( .B(arr[873]), .A(arr[889]), .S(n1100), .Y(n650) );
  MUX2X1 U3200 ( .B(arr[841]), .A(arr[857]), .S(n1100), .Y(n649) );
  MUX2X1 U3201 ( .B(arr[809]), .A(arr[825]), .S(n1100), .Y(n653) );
  MUX2X1 U3202 ( .B(arr[777]), .A(arr[793]), .S(n1100), .Y(n652) );
  MUX2X1 U3203 ( .B(n651), .A(n648), .S(n1183), .Y(n655) );
  MUX2X1 U3204 ( .B(arr[745]), .A(arr[761]), .S(n1101), .Y(n659) );
  MUX2X1 U3205 ( .B(arr[713]), .A(arr[729]), .S(n1101), .Y(n658) );
  MUX2X1 U3206 ( .B(arr[681]), .A(arr[697]), .S(n1101), .Y(n662) );
  MUX2X1 U3207 ( .B(arr[649]), .A(arr[665]), .S(n1101), .Y(n661) );
  MUX2X1 U3208 ( .B(n660), .A(n657), .S(n1183), .Y(n671) );
  MUX2X1 U3209 ( .B(arr[617]), .A(arr[633]), .S(n1101), .Y(n665) );
  MUX2X1 U3210 ( .B(arr[585]), .A(arr[601]), .S(n1101), .Y(n664) );
  MUX2X1 U3211 ( .B(arr[553]), .A(arr[569]), .S(n1101), .Y(n668) );
  MUX2X1 U3212 ( .B(arr[521]), .A(arr[537]), .S(n1101), .Y(n667) );
  MUX2X1 U3213 ( .B(n666), .A(n663), .S(n1183), .Y(n670) );
  MUX2X1 U3214 ( .B(n669), .A(n654), .S(n17), .Y(n703) );
  MUX2X1 U3215 ( .B(arr[489]), .A(arr[505]), .S(n1101), .Y(n674) );
  MUX2X1 U3216 ( .B(arr[457]), .A(arr[473]), .S(n1101), .Y(n673) );
  MUX2X1 U3217 ( .B(arr[425]), .A(arr[441]), .S(n1101), .Y(n677) );
  MUX2X1 U3218 ( .B(arr[393]), .A(arr[409]), .S(n1101), .Y(n676) );
  MUX2X1 U3219 ( .B(n675), .A(n672), .S(n1183), .Y(n686) );
  MUX2X1 U3220 ( .B(arr[361]), .A(arr[377]), .S(n1102), .Y(n680) );
  MUX2X1 U3221 ( .B(arr[329]), .A(arr[345]), .S(n1102), .Y(n679) );
  MUX2X1 U3222 ( .B(arr[297]), .A(arr[313]), .S(n1102), .Y(n683) );
  MUX2X1 U3223 ( .B(arr[265]), .A(arr[281]), .S(n1102), .Y(n682) );
  MUX2X1 U3224 ( .B(n681), .A(n678), .S(n1183), .Y(n685) );
  MUX2X1 U3225 ( .B(arr[233]), .A(arr[249]), .S(n1102), .Y(n689) );
  MUX2X1 U3226 ( .B(arr[201]), .A(arr[217]), .S(n1102), .Y(n688) );
  MUX2X1 U3227 ( .B(arr[169]), .A(arr[185]), .S(n1102), .Y(n692) );
  MUX2X1 U3228 ( .B(arr[137]), .A(arr[153]), .S(n1102), .Y(n691) );
  MUX2X1 U3229 ( .B(n690), .A(n687), .S(n1183), .Y(n701) );
  MUX2X1 U3230 ( .B(arr[105]), .A(arr[121]), .S(n1102), .Y(n695) );
  MUX2X1 U3231 ( .B(arr[73]), .A(arr[89]), .S(n1102), .Y(n694) );
  MUX2X1 U3232 ( .B(arr[41]), .A(arr[57]), .S(n1102), .Y(n698) );
  MUX2X1 U3233 ( .B(arr[9]), .A(arr[25]), .S(n1102), .Y(n697) );
  MUX2X1 U3234 ( .B(n696), .A(n693), .S(n1183), .Y(n700) );
  MUX2X1 U3235 ( .B(n699), .A(n684), .S(n17), .Y(n702) );
  MUX2X1 U3236 ( .B(arr[1002]), .A(arr[1018]), .S(n1103), .Y(n706) );
  MUX2X1 U3237 ( .B(arr[970]), .A(arr[986]), .S(n1103), .Y(n705) );
  MUX2X1 U3238 ( .B(arr[938]), .A(arr[954]), .S(n1103), .Y(n709) );
  MUX2X1 U3239 ( .B(arr[906]), .A(arr[922]), .S(n1103), .Y(n708) );
  MUX2X1 U3240 ( .B(n707), .A(n704), .S(n1184), .Y(n718) );
  MUX2X1 U3241 ( .B(arr[874]), .A(arr[890]), .S(n1103), .Y(n712) );
  MUX2X1 U3242 ( .B(arr[842]), .A(arr[858]), .S(n1103), .Y(n711) );
  MUX2X1 U3243 ( .B(arr[810]), .A(arr[826]), .S(n1103), .Y(n715) );
  MUX2X1 U3244 ( .B(arr[778]), .A(arr[794]), .S(n1103), .Y(n714) );
  MUX2X1 U3245 ( .B(n713), .A(n710), .S(n1184), .Y(n717) );
  MUX2X1 U3246 ( .B(arr[746]), .A(arr[762]), .S(n1103), .Y(n721) );
  MUX2X1 U3247 ( .B(arr[714]), .A(arr[730]), .S(n1103), .Y(n720) );
  MUX2X1 U3248 ( .B(arr[682]), .A(arr[698]), .S(n1103), .Y(n724) );
  MUX2X1 U3249 ( .B(arr[650]), .A(arr[666]), .S(n1103), .Y(n723) );
  MUX2X1 U3250 ( .B(n722), .A(n719), .S(n1184), .Y(n733) );
  MUX2X1 U3251 ( .B(arr[618]), .A(arr[634]), .S(n1104), .Y(n727) );
  MUX2X1 U3252 ( .B(arr[586]), .A(arr[602]), .S(n1104), .Y(n726) );
  MUX2X1 U3253 ( .B(arr[554]), .A(arr[570]), .S(n1104), .Y(n730) );
  MUX2X1 U3254 ( .B(arr[522]), .A(arr[538]), .S(n1104), .Y(n729) );
  MUX2X1 U3255 ( .B(n728), .A(n725), .S(n1184), .Y(n732) );
  MUX2X1 U3256 ( .B(n731), .A(n716), .S(n17), .Y(n765) );
  MUX2X1 U3257 ( .B(arr[490]), .A(arr[506]), .S(n1104), .Y(n736) );
  MUX2X1 U3258 ( .B(arr[458]), .A(arr[474]), .S(n1104), .Y(n735) );
  MUX2X1 U3259 ( .B(arr[426]), .A(arr[442]), .S(n1104), .Y(n739) );
  MUX2X1 U3260 ( .B(arr[394]), .A(arr[410]), .S(n1104), .Y(n738) );
  MUX2X1 U3261 ( .B(n737), .A(n734), .S(n1184), .Y(n748) );
  MUX2X1 U3262 ( .B(arr[362]), .A(arr[378]), .S(n1104), .Y(n742) );
  MUX2X1 U3263 ( .B(arr[330]), .A(arr[346]), .S(n1104), .Y(n741) );
  MUX2X1 U3264 ( .B(arr[298]), .A(arr[314]), .S(n1104), .Y(n745) );
  MUX2X1 U3265 ( .B(arr[266]), .A(arr[282]), .S(n1104), .Y(n744) );
  MUX2X1 U3266 ( .B(n743), .A(n740), .S(n1184), .Y(n747) );
  MUX2X1 U3267 ( .B(arr[234]), .A(arr[250]), .S(n1105), .Y(n751) );
  MUX2X1 U3268 ( .B(arr[202]), .A(arr[218]), .S(n1105), .Y(n750) );
  MUX2X1 U3269 ( .B(arr[170]), .A(arr[186]), .S(n1105), .Y(n754) );
  MUX2X1 U3270 ( .B(arr[138]), .A(arr[154]), .S(n1105), .Y(n753) );
  MUX2X1 U3271 ( .B(n752), .A(n749), .S(n1184), .Y(n763) );
  MUX2X1 U3272 ( .B(arr[106]), .A(arr[122]), .S(n1105), .Y(n757) );
  MUX2X1 U3273 ( .B(arr[74]), .A(arr[90]), .S(n1105), .Y(n756) );
  MUX2X1 U3274 ( .B(arr[42]), .A(arr[58]), .S(n1105), .Y(n760) );
  MUX2X1 U3275 ( .B(arr[10]), .A(arr[26]), .S(n1105), .Y(n759) );
  MUX2X1 U3276 ( .B(n758), .A(n755), .S(n1184), .Y(n762) );
  MUX2X1 U3277 ( .B(n761), .A(n746), .S(n17), .Y(n764) );
  MUX2X1 U3278 ( .B(arr[1003]), .A(arr[1019]), .S(n1105), .Y(n768) );
  MUX2X1 U3279 ( .B(arr[971]), .A(arr[987]), .S(n1105), .Y(n767) );
  MUX2X1 U3280 ( .B(arr[939]), .A(arr[955]), .S(n1105), .Y(n771) );
  MUX2X1 U3281 ( .B(arr[907]), .A(arr[923]), .S(n1105), .Y(n770) );
  MUX2X1 U3282 ( .B(n769), .A(n766), .S(n1184), .Y(n780) );
  MUX2X1 U3283 ( .B(arr[875]), .A(arr[891]), .S(n1106), .Y(n774) );
  MUX2X1 U3284 ( .B(arr[843]), .A(arr[859]), .S(n1106), .Y(n773) );
  MUX2X1 U3285 ( .B(arr[811]), .A(arr[827]), .S(n1106), .Y(n777) );
  MUX2X1 U3286 ( .B(arr[779]), .A(arr[795]), .S(n1106), .Y(n776) );
  MUX2X1 U3287 ( .B(n775), .A(n772), .S(n1184), .Y(n779) );
  MUX2X1 U3288 ( .B(arr[747]), .A(arr[763]), .S(n1106), .Y(n783) );
  MUX2X1 U3289 ( .B(arr[715]), .A(arr[731]), .S(n1106), .Y(n782) );
  MUX2X1 U3290 ( .B(arr[683]), .A(arr[699]), .S(n1106), .Y(n786) );
  MUX2X1 U3291 ( .B(arr[651]), .A(arr[667]), .S(n1106), .Y(n785) );
  MUX2X1 U3292 ( .B(n784), .A(n781), .S(n1184), .Y(n795) );
  MUX2X1 U3293 ( .B(arr[619]), .A(arr[635]), .S(n1106), .Y(n789) );
  MUX2X1 U3294 ( .B(arr[587]), .A(arr[603]), .S(n1106), .Y(n788) );
  MUX2X1 U3295 ( .B(arr[555]), .A(arr[571]), .S(n1106), .Y(n792) );
  MUX2X1 U3296 ( .B(arr[523]), .A(arr[539]), .S(n1106), .Y(n791) );
  MUX2X1 U3297 ( .B(n790), .A(n787), .S(n1184), .Y(n794) );
  MUX2X1 U3298 ( .B(n793), .A(n778), .S(n17), .Y(n827) );
  MUX2X1 U3299 ( .B(arr[491]), .A(arr[507]), .S(n1107), .Y(n798) );
  MUX2X1 U3300 ( .B(arr[459]), .A(arr[475]), .S(n1107), .Y(n797) );
  MUX2X1 U3301 ( .B(arr[427]), .A(arr[443]), .S(n1107), .Y(n801) );
  MUX2X1 U3302 ( .B(arr[395]), .A(arr[411]), .S(n1107), .Y(n800) );
  MUX2X1 U3303 ( .B(n799), .A(n796), .S(n1185), .Y(n810) );
  MUX2X1 U3304 ( .B(arr[363]), .A(arr[379]), .S(n1107), .Y(n804) );
  MUX2X1 U3305 ( .B(arr[331]), .A(arr[347]), .S(n1107), .Y(n803) );
  MUX2X1 U3306 ( .B(arr[299]), .A(arr[315]), .S(n1107), .Y(n807) );
  MUX2X1 U3307 ( .B(arr[267]), .A(arr[283]), .S(n1107), .Y(n806) );
  MUX2X1 U3308 ( .B(n805), .A(n802), .S(n1185), .Y(n809) );
  MUX2X1 U3309 ( .B(arr[235]), .A(arr[251]), .S(n1107), .Y(n813) );
  MUX2X1 U3310 ( .B(arr[203]), .A(arr[219]), .S(n1107), .Y(n812) );
  MUX2X1 U3311 ( .B(arr[171]), .A(arr[187]), .S(n1107), .Y(n816) );
  MUX2X1 U3312 ( .B(arr[139]), .A(arr[155]), .S(n1107), .Y(n815) );
  MUX2X1 U3313 ( .B(n814), .A(n811), .S(n1185), .Y(n825) );
  MUX2X1 U3314 ( .B(arr[107]), .A(arr[123]), .S(n1108), .Y(n819) );
  MUX2X1 U3315 ( .B(arr[75]), .A(arr[91]), .S(n1108), .Y(n818) );
  MUX2X1 U3316 ( .B(arr[43]), .A(arr[59]), .S(n1108), .Y(n822) );
  MUX2X1 U3317 ( .B(arr[11]), .A(arr[27]), .S(n1108), .Y(n821) );
  MUX2X1 U3318 ( .B(n820), .A(n817), .S(n1185), .Y(n824) );
  MUX2X1 U3319 ( .B(n823), .A(n808), .S(n17), .Y(n826) );
  MUX2X1 U3320 ( .B(arr[1004]), .A(arr[1020]), .S(n1108), .Y(n830) );
  MUX2X1 U3321 ( .B(arr[972]), .A(arr[988]), .S(n1108), .Y(n829) );
  MUX2X1 U3322 ( .B(arr[940]), .A(arr[956]), .S(n1108), .Y(n833) );
  MUX2X1 U3323 ( .B(arr[908]), .A(arr[924]), .S(n1108), .Y(n832) );
  MUX2X1 U3324 ( .B(n831), .A(n828), .S(n1185), .Y(n842) );
  MUX2X1 U3325 ( .B(arr[876]), .A(arr[892]), .S(n1108), .Y(n836) );
  MUX2X1 U3326 ( .B(arr[844]), .A(arr[860]), .S(n1108), .Y(n835) );
  MUX2X1 U3327 ( .B(arr[812]), .A(arr[828]), .S(n1108), .Y(n839) );
  MUX2X1 U3328 ( .B(arr[780]), .A(arr[796]), .S(n1108), .Y(n838) );
  MUX2X1 U3329 ( .B(n837), .A(n834), .S(n1185), .Y(n841) );
  MUX2X1 U3330 ( .B(arr[748]), .A(arr[764]), .S(n1109), .Y(n845) );
  MUX2X1 U3331 ( .B(arr[716]), .A(arr[732]), .S(n1109), .Y(n844) );
  MUX2X1 U3332 ( .B(arr[684]), .A(arr[700]), .S(n1109), .Y(n848) );
  MUX2X1 U3333 ( .B(arr[652]), .A(arr[668]), .S(n1109), .Y(n847) );
  MUX2X1 U3334 ( .B(n846), .A(n843), .S(n1185), .Y(n857) );
  MUX2X1 U3335 ( .B(arr[620]), .A(arr[636]), .S(n1109), .Y(n851) );
  MUX2X1 U3336 ( .B(arr[588]), .A(arr[604]), .S(n1109), .Y(n850) );
  MUX2X1 U3337 ( .B(arr[556]), .A(arr[572]), .S(n1109), .Y(n854) );
  MUX2X1 U3338 ( .B(arr[524]), .A(arr[540]), .S(n1109), .Y(n853) );
  MUX2X1 U3339 ( .B(n852), .A(n849), .S(n1185), .Y(n856) );
  MUX2X1 U3340 ( .B(n855), .A(n840), .S(n17), .Y(n889) );
  MUX2X1 U3341 ( .B(arr[492]), .A(arr[508]), .S(n1109), .Y(n860) );
  MUX2X1 U3342 ( .B(arr[460]), .A(arr[476]), .S(n1109), .Y(n859) );
  MUX2X1 U3343 ( .B(arr[428]), .A(arr[444]), .S(n1109), .Y(n863) );
  MUX2X1 U3344 ( .B(arr[396]), .A(arr[412]), .S(n1109), .Y(n862) );
  MUX2X1 U3345 ( .B(n861), .A(n858), .S(n1185), .Y(n872) );
  MUX2X1 U3346 ( .B(arr[364]), .A(arr[380]), .S(n1110), .Y(n866) );
  MUX2X1 U3347 ( .B(arr[332]), .A(arr[348]), .S(n1110), .Y(n865) );
  MUX2X1 U3348 ( .B(arr[300]), .A(arr[316]), .S(n1110), .Y(n869) );
  MUX2X1 U3349 ( .B(arr[268]), .A(arr[284]), .S(n1110), .Y(n868) );
  MUX2X1 U3350 ( .B(n867), .A(n864), .S(n1185), .Y(n871) );
  MUX2X1 U3351 ( .B(arr[236]), .A(arr[252]), .S(n1110), .Y(n875) );
  MUX2X1 U3352 ( .B(arr[204]), .A(arr[220]), .S(n1110), .Y(n874) );
  MUX2X1 U3353 ( .B(arr[172]), .A(arr[188]), .S(n1110), .Y(n878) );
  MUX2X1 U3354 ( .B(arr[140]), .A(arr[156]), .S(n1110), .Y(n877) );
  MUX2X1 U3355 ( .B(n876), .A(n873), .S(n1185), .Y(n887) );
  MUX2X1 U3356 ( .B(arr[108]), .A(arr[124]), .S(n1110), .Y(n881) );
  MUX2X1 U3357 ( .B(arr[76]), .A(arr[92]), .S(n1110), .Y(n880) );
  MUX2X1 U3358 ( .B(arr[44]), .A(arr[60]), .S(n1110), .Y(n884) );
  MUX2X1 U3359 ( .B(arr[12]), .A(arr[28]), .S(n1110), .Y(n883) );
  MUX2X1 U3360 ( .B(n882), .A(n879), .S(n1185), .Y(n886) );
  MUX2X1 U3361 ( .B(n885), .A(n870), .S(n17), .Y(n888) );
  MUX2X1 U3362 ( .B(arr[1005]), .A(arr[1021]), .S(n1111), .Y(n892) );
  MUX2X1 U3363 ( .B(arr[973]), .A(arr[989]), .S(n1111), .Y(n891) );
  MUX2X1 U3364 ( .B(arr[941]), .A(arr[957]), .S(n1111), .Y(n895) );
  MUX2X1 U3365 ( .B(arr[909]), .A(arr[925]), .S(n1111), .Y(n894) );
  MUX2X1 U3366 ( .B(n893), .A(n890), .S(n1186), .Y(n904) );
  MUX2X1 U3367 ( .B(arr[877]), .A(arr[893]), .S(n1111), .Y(n898) );
  MUX2X1 U3368 ( .B(arr[845]), .A(arr[861]), .S(n1111), .Y(n897) );
  MUX2X1 U3369 ( .B(arr[813]), .A(arr[829]), .S(n1111), .Y(n901) );
  MUX2X1 U3370 ( .B(arr[781]), .A(arr[797]), .S(n1111), .Y(n900) );
  MUX2X1 U3371 ( .B(n899), .A(n896), .S(n1186), .Y(n903) );
  MUX2X1 U3372 ( .B(arr[749]), .A(arr[765]), .S(n1111), .Y(n907) );
  MUX2X1 U3373 ( .B(arr[717]), .A(arr[733]), .S(n1111), .Y(n906) );
  MUX2X1 U3374 ( .B(arr[685]), .A(arr[701]), .S(n1111), .Y(n910) );
  MUX2X1 U3375 ( .B(arr[653]), .A(arr[669]), .S(n1111), .Y(n909) );
  MUX2X1 U3376 ( .B(n908), .A(n905), .S(n1186), .Y(n919) );
  MUX2X1 U3377 ( .B(arr[621]), .A(arr[637]), .S(n1112), .Y(n913) );
  MUX2X1 U3378 ( .B(arr[589]), .A(arr[605]), .S(n1112), .Y(n912) );
  MUX2X1 U3379 ( .B(arr[557]), .A(arr[573]), .S(n1112), .Y(n916) );
  MUX2X1 U3380 ( .B(arr[525]), .A(arr[541]), .S(n1112), .Y(n915) );
  MUX2X1 U3381 ( .B(n914), .A(n911), .S(n1186), .Y(n918) );
  MUX2X1 U3382 ( .B(n917), .A(n902), .S(n17), .Y(n951) );
  MUX2X1 U3383 ( .B(arr[493]), .A(arr[509]), .S(n1112), .Y(n922) );
  MUX2X1 U3384 ( .B(arr[461]), .A(arr[477]), .S(n1112), .Y(n921) );
  MUX2X1 U3385 ( .B(arr[429]), .A(arr[445]), .S(n1112), .Y(n925) );
  MUX2X1 U3386 ( .B(arr[397]), .A(arr[413]), .S(n1112), .Y(n924) );
  MUX2X1 U3387 ( .B(n923), .A(n920), .S(n1186), .Y(n934) );
  MUX2X1 U3388 ( .B(arr[365]), .A(arr[381]), .S(n1112), .Y(n928) );
  MUX2X1 U3389 ( .B(arr[333]), .A(arr[349]), .S(n1112), .Y(n927) );
  MUX2X1 U3390 ( .B(arr[301]), .A(arr[317]), .S(n1112), .Y(n931) );
  MUX2X1 U3391 ( .B(arr[269]), .A(arr[285]), .S(n1112), .Y(n930) );
  MUX2X1 U3392 ( .B(n929), .A(n926), .S(n1186), .Y(n933) );
  MUX2X1 U3393 ( .B(arr[237]), .A(arr[253]), .S(n1113), .Y(n937) );
  MUX2X1 U3394 ( .B(arr[205]), .A(arr[221]), .S(n1113), .Y(n936) );
  MUX2X1 U3395 ( .B(arr[173]), .A(arr[189]), .S(n1113), .Y(n940) );
  MUX2X1 U3396 ( .B(arr[141]), .A(arr[157]), .S(n1113), .Y(n939) );
  MUX2X1 U3397 ( .B(n938), .A(n935), .S(n1186), .Y(n949) );
  MUX2X1 U3398 ( .B(arr[109]), .A(arr[125]), .S(n1113), .Y(n943) );
  MUX2X1 U3399 ( .B(arr[77]), .A(arr[93]), .S(n1113), .Y(n942) );
  MUX2X1 U3400 ( .B(arr[45]), .A(arr[61]), .S(n1113), .Y(n946) );
  MUX2X1 U3401 ( .B(arr[13]), .A(arr[29]), .S(n1113), .Y(n945) );
  MUX2X1 U3402 ( .B(n944), .A(n941), .S(n1186), .Y(n948) );
  MUX2X1 U3403 ( .B(n947), .A(n932), .S(n17), .Y(n950) );
  MUX2X1 U3404 ( .B(arr[1006]), .A(arr[1022]), .S(n1113), .Y(n954) );
  MUX2X1 U3405 ( .B(arr[974]), .A(arr[990]), .S(n1113), .Y(n953) );
  MUX2X1 U3406 ( .B(arr[942]), .A(arr[958]), .S(n1113), .Y(n957) );
  MUX2X1 U3407 ( .B(arr[910]), .A(arr[926]), .S(n1113), .Y(n956) );
  MUX2X1 U3408 ( .B(n955), .A(n952), .S(n1186), .Y(n966) );
  MUX2X1 U3409 ( .B(arr[878]), .A(arr[894]), .S(n1114), .Y(n960) );
  MUX2X1 U3410 ( .B(arr[846]), .A(arr[862]), .S(n1114), .Y(n959) );
  MUX2X1 U3411 ( .B(arr[814]), .A(arr[830]), .S(n1114), .Y(n963) );
  MUX2X1 U3412 ( .B(arr[782]), .A(arr[798]), .S(n1114), .Y(n962) );
  MUX2X1 U3413 ( .B(n961), .A(n958), .S(n1186), .Y(n965) );
  MUX2X1 U3414 ( .B(arr[750]), .A(arr[766]), .S(n1114), .Y(n969) );
  MUX2X1 U3415 ( .B(arr[718]), .A(arr[734]), .S(n1114), .Y(n968) );
  MUX2X1 U3416 ( .B(arr[686]), .A(arr[702]), .S(n1114), .Y(n972) );
  MUX2X1 U3417 ( .B(arr[654]), .A(arr[670]), .S(n1114), .Y(n971) );
  MUX2X1 U3418 ( .B(n970), .A(n967), .S(n1186), .Y(n981) );
  MUX2X1 U3419 ( .B(arr[622]), .A(arr[638]), .S(n1114), .Y(n975) );
  MUX2X1 U3420 ( .B(arr[590]), .A(arr[606]), .S(n1114), .Y(n974) );
  MUX2X1 U3421 ( .B(arr[558]), .A(arr[574]), .S(n1114), .Y(n978) );
  MUX2X1 U3422 ( .B(arr[526]), .A(arr[542]), .S(n1114), .Y(n977) );
  MUX2X1 U3423 ( .B(n976), .A(n973), .S(n1186), .Y(n980) );
  MUX2X1 U3424 ( .B(n979), .A(n964), .S(n17), .Y(n1013) );
  MUX2X1 U3425 ( .B(arr[494]), .A(arr[510]), .S(n1115), .Y(n984) );
  MUX2X1 U3426 ( .B(arr[462]), .A(arr[478]), .S(n1115), .Y(n983) );
  MUX2X1 U3427 ( .B(arr[430]), .A(arr[446]), .S(n1115), .Y(n987) );
  MUX2X1 U3428 ( .B(arr[398]), .A(arr[414]), .S(n1115), .Y(n986) );
  MUX2X1 U3429 ( .B(n985), .A(n982), .S(n1187), .Y(n996) );
  MUX2X1 U3430 ( .B(arr[366]), .A(arr[382]), .S(n1115), .Y(n990) );
  MUX2X1 U3431 ( .B(arr[334]), .A(arr[350]), .S(n1115), .Y(n989) );
  MUX2X1 U3432 ( .B(arr[302]), .A(arr[318]), .S(n1115), .Y(n993) );
  MUX2X1 U3433 ( .B(arr[270]), .A(arr[286]), .S(n1115), .Y(n992) );
  MUX2X1 U3434 ( .B(n991), .A(n988), .S(n1187), .Y(n995) );
  MUX2X1 U3435 ( .B(arr[238]), .A(arr[254]), .S(n1115), .Y(n999) );
  MUX2X1 U3436 ( .B(arr[206]), .A(arr[222]), .S(n1115), .Y(n998) );
  MUX2X1 U3437 ( .B(arr[174]), .A(arr[190]), .S(n1115), .Y(n1002) );
  MUX2X1 U3438 ( .B(arr[142]), .A(arr[158]), .S(n1115), .Y(n1001) );
  MUX2X1 U3439 ( .B(n1000), .A(n997), .S(n1187), .Y(n1011) );
  MUX2X1 U3440 ( .B(arr[110]), .A(arr[126]), .S(n1116), .Y(n1005) );
  MUX2X1 U3441 ( .B(arr[78]), .A(arr[94]), .S(n1116), .Y(n1004) );
  MUX2X1 U3442 ( .B(arr[46]), .A(arr[62]), .S(n1116), .Y(n1008) );
  MUX2X1 U3443 ( .B(arr[14]), .A(arr[30]), .S(n1116), .Y(n1007) );
  MUX2X1 U3444 ( .B(n1006), .A(n1003), .S(n1187), .Y(n1010) );
  MUX2X1 U3445 ( .B(n1009), .A(n994), .S(n17), .Y(n1012) );
  MUX2X1 U3446 ( .B(arr[1007]), .A(arr[1023]), .S(n1116), .Y(n1016) );
  MUX2X1 U3447 ( .B(arr[975]), .A(arr[991]), .S(n1116), .Y(n1015) );
  MUX2X1 U3448 ( .B(arr[943]), .A(arr[959]), .S(n1116), .Y(n1019) );
  MUX2X1 U3449 ( .B(arr[911]), .A(arr[927]), .S(n1116), .Y(n1018) );
  MUX2X1 U3450 ( .B(n1017), .A(n1014), .S(n1187), .Y(n1028) );
  MUX2X1 U3451 ( .B(arr[879]), .A(arr[895]), .S(n1116), .Y(n1022) );
  MUX2X1 U3452 ( .B(arr[847]), .A(arr[863]), .S(n1116), .Y(n1021) );
  MUX2X1 U3453 ( .B(arr[815]), .A(arr[831]), .S(n1116), .Y(n1025) );
  MUX2X1 U3454 ( .B(arr[783]), .A(arr[799]), .S(n1116), .Y(n1024) );
  MUX2X1 U3455 ( .B(n1023), .A(n1020), .S(n1187), .Y(n1027) );
  MUX2X1 U3456 ( .B(arr[751]), .A(arr[767]), .S(n1117), .Y(n1031) );
  MUX2X1 U3457 ( .B(arr[719]), .A(arr[735]), .S(n1117), .Y(n1030) );
  MUX2X1 U3458 ( .B(arr[687]), .A(arr[703]), .S(n1117), .Y(n1034) );
  MUX2X1 U3459 ( .B(arr[655]), .A(arr[671]), .S(n1117), .Y(n1033) );
  MUX2X1 U3460 ( .B(n1032), .A(n1029), .S(n1187), .Y(n1043) );
  MUX2X1 U3461 ( .B(arr[623]), .A(arr[639]), .S(n1117), .Y(n1037) );
  MUX2X1 U3462 ( .B(arr[591]), .A(arr[607]), .S(n1117), .Y(n1036) );
  MUX2X1 U3463 ( .B(arr[559]), .A(arr[575]), .S(n1117), .Y(n1040) );
  MUX2X1 U3464 ( .B(arr[527]), .A(arr[543]), .S(n1117), .Y(n1039) );
  MUX2X1 U3465 ( .B(n1038), .A(n1035), .S(n1187), .Y(n1042) );
  MUX2X1 U3466 ( .B(n1041), .A(n1026), .S(n17), .Y(n1075) );
  MUX2X1 U3467 ( .B(arr[495]), .A(arr[511]), .S(n1117), .Y(n1046) );
  MUX2X1 U3468 ( .B(arr[463]), .A(arr[479]), .S(n1117), .Y(n1045) );
  MUX2X1 U3469 ( .B(arr[431]), .A(arr[447]), .S(n1117), .Y(n1049) );
  MUX2X1 U3470 ( .B(arr[399]), .A(arr[415]), .S(n1117), .Y(n1048) );
  MUX2X1 U3471 ( .B(n1047), .A(n1044), .S(n1187), .Y(n1058) );
  MUX2X1 U3472 ( .B(arr[367]), .A(arr[383]), .S(n1118), .Y(n1052) );
  MUX2X1 U3473 ( .B(arr[335]), .A(arr[351]), .S(n1118), .Y(n1051) );
  MUX2X1 U3474 ( .B(arr[303]), .A(arr[319]), .S(n1118), .Y(n1055) );
  MUX2X1 U3475 ( .B(arr[271]), .A(arr[287]), .S(n1118), .Y(n1054) );
  MUX2X1 U3476 ( .B(n1053), .A(n1050), .S(n1187), .Y(n1057) );
  MUX2X1 U3477 ( .B(arr[239]), .A(arr[255]), .S(n1118), .Y(n1061) );
  MUX2X1 U3478 ( .B(arr[207]), .A(arr[223]), .S(n1118), .Y(n1060) );
  MUX2X1 U3479 ( .B(arr[175]), .A(arr[191]), .S(n1118), .Y(n1064) );
  MUX2X1 U3480 ( .B(arr[143]), .A(arr[159]), .S(n1118), .Y(n1063) );
  MUX2X1 U3481 ( .B(n1062), .A(n1059), .S(n1187), .Y(n1073) );
  MUX2X1 U3482 ( .B(arr[111]), .A(arr[127]), .S(n1118), .Y(n1067) );
  MUX2X1 U3483 ( .B(arr[79]), .A(arr[95]), .S(n1118), .Y(n1066) );
  MUX2X1 U3484 ( .B(arr[47]), .A(arr[63]), .S(n1118), .Y(n1070) );
  MUX2X1 U3485 ( .B(arr[15]), .A(arr[31]), .S(n1118), .Y(n1069) );
  MUX2X1 U3486 ( .B(n1068), .A(n1065), .S(n1187), .Y(n1072) );
  MUX2X1 U3487 ( .B(n1071), .A(n1056), .S(n17), .Y(n1074) );
  AND2X2 U3488 ( .A(n3440), .B(n3439), .Y(n2870) );
  INVX1 U3489 ( .A(n3440), .Y(n3438) );
  INVX1 U3490 ( .A(fillcount[5]), .Y(n3442) );
  AND2X2 U3491 ( .A(n3413), .B(wr_ptr[0]), .Y(n2907) );
  AND2X2 U3492 ( .A(n3413), .B(n2852), .Y(n2889) );
  AND2X2 U3493 ( .A(wr_ptr[0]), .B(n2851), .Y(n2342) );
  AND2X2 U3494 ( .A(n2851), .B(n2852), .Y(n2323) );
endmodule


module ddr2_controller ( dout, raddr, fillcount, notfull, ready, ck_pad, 
        ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad, webar_pad, 
        ba_pad, a_pad, dm_pad, odt_pad, dq_pad, dqs_pad, dqsbar_pad, clk, 
        reset, read, cmd, din, addr, initddr );
  output [15:0] dout;
  output [24:0] raddr;
  output [6:0] fillcount;
  output [1:0] ba_pad;
  output [12:0] a_pad;
  output [1:0] dm_pad;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] cmd;
  input [15:0] din;
  input [24:0] addr;
  input clk, reset, read, initddr;
  output notfull, ready, ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad,
         casbar_pad, webar_pad, odt_pad;
  wire   ck_i, n7, full, init_rasbar, init_casbar, init_webar, init_odt,
         init_cke, rasbar_i, casbar_i, webar_i, n11, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134;
  wire   [32:0] CMD_data_in;
  wire   [40:0] RETURN_data_in;
  wire   [1:0] init_ba;
  wire   [12:0] init_a;
  wire   [12:0] a_i;
  wire   [1:0] ba_i;
  wire   [15:0] dq_i;
  wire   [1:0] dqs_i;
  wire   [1:0] dqsbar_i;
  wire   [1:0] dm_i;

  DFFPOSX1 ck_i_reg ( .D(n7), .CLK(clk), .Q(ck_i) );
  INVX2 U3 ( .A(full), .Y(notfull) );
  AND2X1 U5 ( .A(init_webar), .B(n11), .Y(webar_i) );
  AND2X1 U6 ( .A(init_rasbar), .B(n11), .Y(rasbar_i) );
  NOR2X1 U7 ( .A(reset), .B(ck_i), .Y(n7) );
  AND2X1 U9 ( .A(init_casbar), .B(n11), .Y(casbar_i) );
  AND2X1 U10 ( .A(init_ba[1]), .B(n11), .Y(ba_i[1]) );
  AND2X1 U11 ( .A(init_ba[0]), .B(n11), .Y(ba_i[0]) );
  AND2X1 U12 ( .A(init_a[9]), .B(n11), .Y(a_i[9]) );
  AND2X1 U13 ( .A(init_a[8]), .B(n11), .Y(a_i[8]) );
  AND2X1 U14 ( .A(init_a[7]), .B(n11), .Y(a_i[7]) );
  AND2X1 U16 ( .A(init_a[5]), .B(n11), .Y(a_i[5]) );
  AND2X1 U17 ( .A(init_a[4]), .B(n11), .Y(a_i[4]) );
  AND2X1 U18 ( .A(init_a[3]), .B(n11), .Y(a_i[3]) );
  AND2X1 U19 ( .A(init_a[2]), .B(n11), .Y(a_i[2]) );
  AND2X1 U20 ( .A(init_a[1]), .B(n11), .Y(a_i[1]) );
  AND2X1 U23 ( .A(init_a[10]), .B(n11), .Y(a_i[10]) );
  AND2X1 U24 ( .A(init_a[0]), .B(n11), .Y(a_i[0]) );
  FIFO_DEPTH_P26_WIDTH16 FIFO_IN ( .clk(clk), .reset(reset), .data_in(din), 
        .put(1'b0), .get(1'b0), .data_out({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16}), .empty(SYNOPSYS_UNCONNECTED_17), .full(full), .fillcount(fillcount) );
  FIFO_DEPTH_P26_WIDTH33 FIFO_CMD ( .clk(clk), .reset(reset), .data_in({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .put(1'b0), .get(
        1'b0), .data_out({SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50}), .empty(SYNOPSYS_UNCONNECTED_51), .full(
        SYNOPSYS_UNCONNECTED_52), .fillcount({SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59}) );
  FIFO_DEPTH_P26_WIDTH41 FIFO_RETURN ( .clk(clk), .reset(reset), .data_in({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .put(1'b0), .get(1'b0), .data_out({
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100}), .empty(SYNOPSYS_UNCONNECTED_101), .full(
        SYNOPSYS_UNCONNECTED_102), .fillcount({SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109}) );
  ddr2_init_engine XINIT ( .ready(ready), .csbar(SYNOPSYS_UNCONNECTED_110), 
        .rasbar(init_rasbar), .casbar(init_casbar), .webar(init_webar), .ba(
        init_ba), .a({SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112, 
        init_a[10:7], SYNOPSYS_UNCONNECTED_113, init_a[5:0]}), .odt(init_odt), 
        .ts_con(SYNOPSYS_UNCONNECTED_114), .cke(init_cke), .clk(clk), .reset(
        reset), .init(initddr), .ck(1'b0) );
  SSTL18DDR2INTERFACE XSSTL ( .ck_pad(ck_pad), .ckbar_pad(ckbar_pad), 
        .cke_pad(cke_pad), .csbar_pad(csbar_pad), .rasbar_pad(rasbar_pad), 
        .casbar_pad(casbar_pad), .webar_pad(webar_pad), .ba_pad(ba_pad), 
        .a_pad(a_pad), .dm_pad(dm_pad), .odt_pad(odt_pad), .dq_o({
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, 
        SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, 
        SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120, 
        SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130}), .dqs_o({
        SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132}), .dqsbar_o({
        SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134}), .dq_pad(dq_pad), 
        .dqs_pad(dqs_pad), .dqsbar_pad(dqsbar_pad), .ri_i(1'b0), .ts_i(1'b0), 
        .ck_i(ck_i), .cke_i(init_cke), .csbar_i(1'b0), .rasbar_i(rasbar_i), 
        .casbar_i(casbar_i), .webar_i(webar_i), .ba_i(ba_i), .a_i({1'b0, 1'b0, 
        a_i[10:7], 1'b0, a_i[5:0]}), .dq_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dqs_i({
        1'b0, 1'b0}), .dqsbar_i({1'b0, 1'b0}), .dm_i({1'b0, 1'b0}), .odt_i(
        init_odt) );
  INVX2 U25 ( .A(ready), .Y(n11) );
endmodule

